* NGSPICE file created from team_10_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt team_10_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3155_ _1564_ _1583_ _0906_ _1562_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2106_ team_10_WB.instance_to_wrap.dispFSM.guesses\[6\] net114 net138 net834 vssd1
+ vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3086_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _1537_ net200 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[79\] sky130_fd_sc_hd__mux2_1
XFILLER_0_89_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2037_ team_10_WB.instance_to_wrap.dispFSM.guesses\[75\] net111 net136 team_10_WB.instance_to_wrap.dispFSM.msg\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3443__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3988_ clknet_leaf_44_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[25\]
+ _0056_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2939_ net210 net150 net121 net810 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[44\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4502__313 vssd1 vssd1 vccd1 vccd1 _4502__313/HI net313 sky130_fd_sc_hd__conb_1
XANTENNA__3286__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2190__A team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2954__B2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4609_ net383 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4663__431 vssd1 vssd1 vccd1 vccd1 _4663__431/HI net431 sky130_fd_sc_hd__conb_1
XFILLER_0_115_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4580__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4704__472 vssd1 vssd1 vccd1 vccd1 _4704__472/HI net472 sky130_fd_sc_hd__conb_1
XFILLER_0_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2275__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3425__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3911_ net243 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3842_ net254 vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3773_ net277 vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2936__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2724_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ _1351_ team_10_WB.instance_to_wrap.clock_div.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _1355_ sky130_fd_sc_hd__a31o_1
XANTENNA__1924__A_N net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2655_ _1308_ _1310_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2586_ _0888_ _0902_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4325_ clknet_leaf_14_wb_clk_i _0715_ _0314_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[48\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_26_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3045__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout127 _1188_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
Xfanout149 net153 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_4
X_4256_ clknet_leaf_56_wb_clk_i _0650_ _0245_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.green
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3113__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3207_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] _1621_ vssd1 vssd1 vccd1
+ vccd1 _1622_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4187_ clknet_leaf_24_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[49\]
+ _0176_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[49\] sky130_fd_sc_hd__dfrtp_1
X_3138_ _1549_ _1567_ _1568_ _1551_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1
+ vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__o32a_1
X_4647__415 vssd1 vssd1 vccd1 vccd1 _4647__415/HI net415 sky130_fd_sc_hd__conb_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2185__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3069_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__mux2_1
XANTENNA__3416__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1978__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4080__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold170 team_10_WB.instance_to_wrap.dispFSM.guesses\[63\] vssd1 vssd1 vccd1 vccd1
+ net722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1
+ net733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\] vssd1 vssd1 vccd1
+ vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2794__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4575__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3407__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2440_ net606 net130 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\]
+ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3343__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2371_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] _1084_ _1144_
+ _1145_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4110_ clknet_leaf_28_wb_clk_i net594 _0109_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4041_ clknet_leaf_31_wb_clk_i net620 _0082_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1902__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3825_ net259 vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2452__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout125_A _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3756_ net292 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2707_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[2\] vssd1 vssd1 vccd1 vccd1 _1345_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3687_ net252 vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2638_ _0922_ _0925_ _0935_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] _0975_
+ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__o221a_1
XFILLER_0_80_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2569_ net220 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] net224 vssd1
+ vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__and3_1
XANTENNA__2252__A_N team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4308_ clknet_leaf_29_wb_clk_i net704 _0297_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4239_ clknet_leaf_50_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[3\]
+ _0228_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1940_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] net144 vssd1 vssd1 vccd1
+ vccd1 _0863_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3261__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1871_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] vssd1 vssd1 vccd1 vccd1
+ _0796_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3610_ net264 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__inv_2
X_4590_ net549 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_0_126_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3541_ net239 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3472_ team_10_WB.instance_to_wrap.dispFSM.guesses\[79\] _1715_ _1842_ _0821_ vssd1
+ vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2423_ net559 _1184_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2354_ _1126_ _1128_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2285_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _1063_ _1064_ _1066_ vssd1
+ vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4024_ clknet_leaf_49_wb_clk_i net611 _0071_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2447__B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout242_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3808_ net281 vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3739_ net278 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2070_ team_10_WB.instance_to_wrap.dispFSM.guesses\[42\] net110 net135 net811 vssd1
+ vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3482__B1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2037__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2972_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] _0835_ net159 vssd1 vssd1 vccd1
+ vccd1 _1487_ sky130_fd_sc_hd__a41o_1
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4711_ net479 vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_0_56_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1923_ net4 net5 net299 vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_17_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4642_ net410 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4573_ net544 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3524_ net238 vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3455_ team_10_WB.instance_to_wrap.host_row2\[54\] net168 net165 team_10_WB.instance_to_wrap.host_row2\[78\]
+ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3842__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2406_ team_10_WB.instance_to_wrap.clock_div.count\[19\] team_10_WB.instance_to_wrap.clock_div.count\[18\]
+ team_10_WB.instance_to_wrap.clock_div.count\[21\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3386_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] net167 net177 team_10_WB.instance_to_wrap.dispFSM.guesses\[43\]
+ _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2337_ _0809_ _0866_ _1093_ _0811_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__a22oi_1
XANTENNA__3053__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2268_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0800_ net211 _0792_ vssd1
+ vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_1286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4007_ clknet_leaf_38_wb_clk_i _0495_ net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2199_ _0984_ _0987_ _0975_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2640__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold30 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] vssd1 vssd1 vccd1 vccd1 net582
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_10_WB.instance_to_wrap.host_row1\[45\] vssd1 vssd1 vccd1 vccd1 net593
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 team_10_WB.instance_to_wrap.host_row1\[63\] vssd1 vssd1 vccd1 vccd1 net604
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 team_10_WB.instance_to_wrap.host_row1\[44\] vssd1 vssd1 vccd1 vccd1 net615
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] vssd1 vssd1 vccd1 vccd1
+ net637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold96 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] vssd1 vssd1 vccd1
+ vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input18_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_5 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3240_ net587 _1642_ net170 vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3171_ _1550_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2122_ net215 net214 team_10_WB.instance_to_wrap.gamelogic.state\[2\] team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__or4b_2
XFILLER_0_59_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2053_ team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] net111 net136 net752 vssd1
+ vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__o22a_1
XANTENNA__2258__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3455__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2258__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4680__448 vssd1 vssd1 vccd1 vccd1 _4680__448/HI net448 sky130_fd_sc_hd__conb_1
XFILLER_0_119_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2955_ _0798_ _1478_ net156 net857 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[7\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1906_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _0829_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4721__489 vssd1 vssd1 vccd1 vccd1 _4721__489/HI net489 sky130_fd_sc_hd__conb_1
XFILLER_0_5_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2886_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] net1 _1467_ vssd1 vssd1 vccd1
+ vccd1 _1468_ sky130_fd_sc_hd__mux2_1
X_4625_ team_10_WB.instance_to_wrap.lcdPlayer.lcd_en vssd1 vssd1 vccd1 vccd1 net77
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4556_ net367 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_114_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout205_A team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2194__B1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3507_ net235 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4487_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[44\]
+ _0470_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3438_ _1719_ _1801_ _1810_ net177 vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3369_ team_10_WB.instance_to_wrap.host_row1\[50\] _1699_ net165 team_10_WB.instance_to_wrap.host_row2\[74\]
+ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2249__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3446__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3382__C1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_102_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2740_ team_10_WB.instance_to_wrap.clock_div.count\[13\] team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ team_10_WB.instance_to_wrap.clock_div.count\[15\] _1362_ vssd1 vssd1 vccd1 vccd1
+ _1365_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2671_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] _1324_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4410_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[7\]
+ _0393_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4341_ clknet_leaf_14_wb_clk_i _0731_ _0330_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[64\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_61_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4272_ clknet_leaf_22_wb_clk_i _0662_ _0261_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3223_ net170 _1631_ _1632_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__nor3_1
XFILLER_0_103_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3154_ net216 _0899_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2105_ team_10_WB.instance_to_wrap.dispFSM.guesses\[15\] net142 net108 net577 vssd1
+ vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a22o_1
X_3085_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__mux2_1
XANTENNA__3428__B1 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2036_ team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] net112 net140 team_10_WB.instance_to_wrap.dispFSM.msg\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3987_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[24\]
+ _0055_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2938_ net211 net150 net121 net804 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[43\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4541__352 vssd1 vssd1 vccd1 vccd1 _4541__352/HI net352 sky130_fd_sc_hd__conb_1
XFILLER_0_60_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2190__B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2869_ team_10_WB.instance_to_wrap.host_message_reg.Cstate net158 _1302_ vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.next_state sky130_fd_sc_hd__a21o_1
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4608_ net382 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4539_ net350 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_130_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3355__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3370__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3910_ net248 vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3841_ net254 vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4525__336 vssd1 vssd1 vccd1 vccd1 _4525__336/HI net336 sky130_fd_sc_hd__conb_1
XFILLER_0_55_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2291__A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3772_ net292 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2723_ net827 _1354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[8\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2654_ _1228_ _1309_ _1315_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_30_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2585_ _1265_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4324_ clknet_leaf_31_wb_clk_i net700 _0313_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3361__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout117 _0875_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout128 _1184_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_4
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_2
X_4255_ clknet_leaf_55_wb_clk_i _0649_ _0244_ vssd1 vssd1 vccd1 vccd1 team_10_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__3850__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3206_ _1621_ _1611_ _1620_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__and3b_1
X_4186_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[48\]
+ _0175_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[48\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4612__386 vssd1 vssd1 vccd1 vccd1 _4612__386/HI net386 sky130_fd_sc_hd__conb_1
X_3137_ _1275_ _1550_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3061__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4686__454 vssd1 vssd1 vccd1 vccd1 _4686__454/HI net454 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3068_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] _1528_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[70\] sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2019_ _0890_ net224 net219 vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4727__495 vssd1 vssd1 vccd1 vccd1 _4727__495/HI net495 sky130_fd_sc_hd__conb_1
XFILLER_0_93_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2388__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold160 team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] vssd1 vssd1 vccd1 vccd1
+ net712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _0730_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3352__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 team_10_WB.instance_to_wrap.host_row1\[60\] vssd1 vssd1 vccd1 vccd1 net734
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold193 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\] vssd1 vssd1 vccd1 vccd1
+ net745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2091__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3343__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2370_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3670__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4040_ clknet_leaf_34_wb_clk_i _0525_ _0081_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3824_ net262 vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2909__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3755_ net272 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2706_ net724 net668 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3686_ net234 vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout118_A _0875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2637_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _1085_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ _1303_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3056__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2568_ _0974_ _1253_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4307_ clknet_leaf_13_wb_clk_i _0697_ _0296_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[30\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2499_ net217 _1218_ _1217_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4238_ clknet_leaf_50_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[2\]
+ _0227_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3098__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4169_ clknet_leaf_46_wb_clk_i _0638_ _0158_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_74_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3325__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4586__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1870_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] vssd1 vssd1 vccd1 vccd1
+ _0795_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3540_ net239 vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3471_ team_10_WB.instance_to_wrap.dispFSM.guesses\[63\] net171 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[15\]
+ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2422_ net156 net155 vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2353_ _1099_ _1124_ _1125_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2284_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _1065_ vssd1 vssd1 vccd1
+ vccd1 _1066_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4023_ clknet_leaf_50_wb_clk_i net562 _0070_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3807_ net279 vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1999_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] net145 net116
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1 vccd1 vccd1 _0750_
+ sky130_fd_sc_hd__o22a_1
X_4787_ net182 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3738_ net290 vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3669_ net287 vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4742__510 vssd1 vssd1 vccd1 vccd1 _4742__510/HI net510 sky130_fd_sc_hd__conb_1
XFILLER_0_112_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4226__534 vssd1 vssd1 vccd1 vccd1 net534 _4226__534/LO sky130_fd_sc_hd__conb_1
XFILLER_0_108_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3467__D1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4093__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2037__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2971_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\] _0834_ net163 vssd1 vssd1 vccd1
+ vccd1 _1486_ sky130_fd_sc_hd__a41o_1
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4710_ net478 vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
XFILLER_0_16_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1922_ net299 net5 vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4641_ net409 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_126_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4572_ net543 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3523_ net230 vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3454_ team_10_WB.instance_to_wrap.host_row1\[70\] _1703_ net177 team_10_WB.instance_to_wrap.host_row2\[70\]
+ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2405_ team_10_WB.instance_to_wrap.clock_div.count\[14\] team_10_WB.instance_to_wrap.clock_div.count\[17\]
+ team_10_WB.instance_to_wrap.clock_div.count\[16\] team_10_WB.instance_to_wrap.clock_div.count\[15\]
+ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3385_ team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] net169 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2336_ _1103_ _1104_ _1105_ _1106_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__and4_1
XANTENNA__2458__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2267_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] _0801_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout185_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4006_ clknet_leaf_41_wb_clk_i _0494_ net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2276__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2198_ _0976_ _0977_ _0980_ _0985_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2433__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold20 team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] vssd1 vssd1 vccd1 vccd1 net572
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _0506_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0581_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1
+ net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_10_WB.instance_to_wrap.host_row1\[47\] vssd1 vssd1 vccd1 vccd1 net616
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] vssd1 vssd1 vccd1
+ vccd1 net627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _0629_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3953__CLK clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_6 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3943__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _0903_ _1277_ _0885_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__and3b_1
XFILLER_0_98_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2121_ team_10_WB.instance_to_wrap.gamelogic.state\[2\] _0923_ team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__and3b_1
XFILLER_0_98_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2052_ team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] net112 net140 net801 vssd1
+ vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__o22a_1
XANTENNA__2258__A2 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2954_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\] net160 _1478_ net209 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[6\] sky130_fd_sc_hd__o22a_1
XFILLER_0_85_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1905_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _0828_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2885_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] net221 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4624_ net393 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4555_ net366 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3391__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3506_ net235 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4486_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[43\]
+ _0469_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_106_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3437_ _1799_ _1803_ _1808_ _1811_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__or4_1
X_3368_ net65 net176 _1746_ net227 vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__o211a_1
XANTENNA__2188__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _0867_ _1090_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3299_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_101_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3134__B1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input30_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4594__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1999__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2948__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2670_ _1324_ _1325_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3373__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4340_ clknet_leaf_31_wb_clk_i net723 _0329_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1923__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4271_ clknet_leaf_49_wb_clk_i _0661_ _0260_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3222_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ _1628_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2479__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3153_ net218 net219 net225 vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2104_ team_10_WB.instance_to_wrap.dispFSM.guesses\[8\] net114 net139 net831 vssd1
+ vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3084_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] _1536_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[78\] sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2035_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] net141 net107 net763 vssd1 vssd1
+ vccd1 vccd1 _0744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3986_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[23\]
+ _0054_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2939__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2937_ net212 net150 net121 net819 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[42\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3059__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2868_ net595 _1455_ _1440_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4607_ net381 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2799_ _1407_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__inv_2
Xhold320 team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\] vssd1 vssd1 vccd1 vccd1
+ net872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4538_ net349 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4469_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[26\]
+ _0452_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4154__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2572__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3840_ net256 vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3310__D_N net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3771_ net271 vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2722_ _1180_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[7\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_89_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2653_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] _0827_ _1225_ _1233_
+ _1313_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__o221a_1
XFILLER_0_120_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2584_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4323_ clknet_leaf_12_wb_clk_i _0713_ _0312_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[46\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_61_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout107 _0915_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout118 _0875_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout129 net130 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4254_ clknet_leaf_51_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[10\]
+ _0243_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3205_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] _1392_ vssd1 vssd1 vccd1 vccd1
+ _1621_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4185_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[47\]
+ _0174_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[47\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3136_ _0903_ _1566_ _1280_ _1277_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3067_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2018_ _0892_ net229 net2 vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__or3b_1
XFILLER_0_89_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2085__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3969_ clknet_leaf_43_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[6\]
+ _0037_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold150 team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] vssd1 vssd1 vccd1
+ vccd1 net702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold161 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\] vssd1 vssd1 vccd1
+ vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold172 team_10_WB.instance_to_wrap.clock_div.count\[1\] vssd1 vssd1 vccd1 vccd1
+ net724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\] vssd1 vssd1 vccd1
+ vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] vssd1 vssd1 vccd1 vccd1
+ net746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4548__359 vssd1 vssd1 vccd1 vccd1 _4548__359/HI net359 sky130_fd_sc_hd__conb_1
XFILLER_0_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3488__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3427__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3823_ net248 vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__inv_2
XANTENNA__3016__C1 team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3754_ net292 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2705_ net668 _1171_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[0\]
+ sky130_fd_sc_hd__nor2_1
X_3685_ net234 vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2636_ net164 _1301_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4653__421 vssd1 vssd1 vccd1 vccd1 _4653__421/HI net421 sky130_fd_sc_hd__conb_1
XFILLER_0_11_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2567_ _1047_ _1252_ net860 vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4306_ clknet_leaf_32_wb_clk_i _0696_ _0295_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2498_ _0812_ _0888_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4237_ clknet_leaf_49_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[1\]
+ _0226_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3072__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4168_ clknet_leaf_46_wb_clk_i _0637_ _0157_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_65_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3119_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1278_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__and3b_1
X_4099_ clknet_leaf_8_wb_clk_i _0570_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3022__A2 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3011__A team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4637__405 vssd1 vssd1 vccd1 vccd1 _4637__405/HI net405 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3470_ team_10_WB.instance_to_wrap.dispFSM.guesses\[23\] net173 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2421_ net163 net153 vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2352_ _1117_ _1122_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2283_ team_10_WB.instance_to_wrap.gamelogic.rights\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4022_ clknet_leaf_50_wb_clk_i net569 _0069_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3806_ net289 vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout130_A _1183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4786_ net533 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XANTENNA_fanout228_A _0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1998_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] net148 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1 vccd1 _0751_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3737_ net289 vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__inv_2
XANTENNA__3067__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3668_ net241 vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2619_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3599_ net285 vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2451__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout290 net296 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2970_ _0835_ net163 vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1921_ net299 net4 vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2442__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ net408 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__2993__B2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4571_ net542 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3522_ net230 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3453_ team_10_WB.instance_to_wrap.host_row2\[86\] _1686_ _1695_ net303 vssd1 vssd1
+ vccd1 vccd1 _1827_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2404_ _1165_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3384_ net66 net175 _1761_ net227 vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2335_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\] _1089_ vssd1 vssd1
+ vccd1 vccd1 _1111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2266_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] net213 vssd1 vssd1 vccd1
+ vccd1 _1048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4005_ clknet_leaf_41_wb_clk_i _0493_ net244 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2197_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] net208 vssd1 vssd1 vccd1
+ vccd1 _0986_ sky130_fd_sc_hd__xor2_1
XANTENNA__3473__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2433__B1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4769_ net180 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3161__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold10 _0508_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 _0511_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_10_WB.instance_to_wrap.clock_div.count\[6\] vssd1 vssd1 vccd1 vccd1 net584
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\] vssd1 vssd1 vccd1
+ vccd1 net595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_10_WB.instance_to_wrap.host_row1\[73\] vssd1 vssd1 vccd1 vccd1 net606
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _0583_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_10_WB.instance_to_wrap.host_row1\[79\] vssd1 vssd1 vccd1 vccd1 net628
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold87 team_10_WB.instance_to_wrap.host_row1\[77\] vssd1 vssd1 vccd1 vccd1 net639
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold98 team_10_WB.instance_to_wrap.host_row1\[65\] vssd1 vssd1 vccd1 vccd1 net650
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2975__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3435__S net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4060__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_4749__517 vssd1 vssd1 vccd1 vccd1 _4749__517/HI net517 sky130_fd_sc_hd__conb_1
X_2120_ net215 net214 vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2051_ team_10_WB.instance_to_wrap.dispFSM.guesses\[69\] net141 net107 net689 vssd1
+ vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3455__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2953_ _0800_ _1478_ _1474_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[5\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1904_ net256 vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2884_ _1222_ _1466_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[4\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_72_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4623_ team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs vssd1 vssd1 vccd1 vccd1 net76
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4554_ net365 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3505_ net236 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4485_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[42\]
+ _0468_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3436_ _1715_ _1720_ net229 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1
+ vccd1 vccd1 _1811_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3367_ net177 _1744_ _1745_ _1743_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout295_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2318_ team_10_WB.instance_to_wrap.host_col\[3\] _0868_ _1092_ net226 _0856_ vssd1
+ vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o311ai_1
XFILLER_0_57_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3298_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2249_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] _0799_ net210 _0794_ _1030_
+ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__a221o_1
XANTENNA__3446__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3382__B2 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_43_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input23_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4564__535 vssd1 vssd1 vccd1 vccd1 net535 _4564__535/LO sky130_fd_sc_hd__conb_1
XFILLER_0_131_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3070__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2948__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1923__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4270_ clknet_leaf_49_wb_clk_i _0660_ _0259_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3221_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ net803 vssd1
+ vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4785__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3152_ team_10_WB.instance_to_wrap.dispFSM.msg\[2\] _1290_ _1550_ _1283_ vssd1 vssd1
+ vccd1 vccd1 _1581_ sky130_fd_sc_hd__o31a_1
XANTENNA__1921__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2103_ team_10_WB.instance_to_wrap.dispFSM.guesses\[9\] net109 net135 net791 vssd1
+ vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__o22a_1
X_3083_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2034_ team_10_WB.instance_to_wrap.dispFSM.guesses\[78\] net113 net137 net740 vssd1
+ vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2100__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3985_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[22\]
+ _0053_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2939__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2936_ net213 net149 net120 net765 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[41\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2867_ _1455_ _1456_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4606_ net380 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2798_ _0815_ net175 _1406_ net293 vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__a211o_2
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold310 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1
+ net862 sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ net348 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xhold321 team_10_WB.instance_to_wrap.clock_div.count\[11\] vssd1 vssd1 vccd1 vccd1
+ net873 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3075__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4468_ clknet_leaf_48_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[25\]
+ _0451_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3116__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3419_ team_10_WB.instance_to_wrap.host_row2\[68\] team_10_WB.instance_to_wrap.dispFSM.guesses\[44\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4399_ clknet_leaf_1_wb_clk_i _0784_ _0382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3104__A team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3052__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4670__438 vssd1 vssd1 vccd1 vccd1 _4670__438/HI net438 sky130_fd_sc_hd__conb_1
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4711__479 vssd1 vssd1 vccd1 vccd1 _4711__479/HI net479 sky130_fd_sc_hd__conb_1
XFILLER_0_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3043__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3770_ net293 vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__inv_2
X_2721_ team_10_WB.instance_to_wrap.clock_div.count\[7\] _1351_ vssd1 vssd1 vccd1
+ vccd1 _1354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2652_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2583_ _1256_ _1258_ _1266_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__or4_1
XFILLER_0_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4322_ clknet_leaf_27_wb_clk_i net674 _0311_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout108 _0915_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
Xfanout119 _0875_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dlymetal6s2s_1
X_4253_ clknet_leaf_51_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[9\]
+ _0242_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3204_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\] _1619_ vssd1 vssd1 vccd1
+ vccd1 _1620_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4184_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[46\]
+ _0173_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[46\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3135_ _1561_ _1565_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3066_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _1527_ net200 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[69\] sky130_fd_sc_hd__mux2_1
XFILLER_0_89_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2017_ net2 net300 _0893_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__2482__B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3034__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3968_ clknet_leaf_43_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[5\]
+ _0036_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2919_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\] net149 net120 net822
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[24\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3899_ net270 vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2702__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold140 team_10_WB.instance_to_wrap.clock_div.count\[13\] vssd1 vssd1 vccd1 vccd1
+ net692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 team_10_WB.instance_to_wrap.dispFSM.guesses\[31\] vssd1 vssd1 vccd1 vccd1
+ net703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold162 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\] vssd1 vssd1 vccd1
+ vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\] vssd1 vssd1 vccd1
+ vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold184 team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] vssd1 vssd1 vccd1 vccd1
+ net736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_10_WB.instance_to_wrap.dispFSM.guesses\[71\] vssd1 vssd1 vccd1 vccd1
+ net747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3949__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2000__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4531__342 vssd1 vssd1 vccd1 vccd1 _4531__342/HI net342 sky130_fd_sc_hd__conb_1
XFILLER_0_95_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3679__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3822_ net259 vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3753_ net284 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2704_ team_10_WB.instance_to_wrap.host_col\[3\] net216 net299 vssd1 vssd1 vccd1
+ vccd1 net81 sky130_fd_sc_hd__mux2_1
XFILLER_0_125_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3684_ net239 vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2635_ _0841_ _1086_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__nor2_2
XFILLER_0_112_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4692__460 vssd1 vssd1 vccd1 vccd1 _4692__460/HI net460 sky130_fd_sc_hd__conb_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2566_ net214 _0948_ net133 vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4305_ clknet_leaf_12_wb_clk_i _0695_ _0294_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2497_ net216 _0891_ _1217_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4236_ clknet_leaf_50_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[0\]
+ _0225_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3098__A3 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4167_ clknet_leaf_46_wb_clk_i _0636_ _0156_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_3118_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] _1278_ vssd1 vssd1 vccd1 vccd1
+ _1549_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4098_ clknet_leaf_8_wb_clk_i _0569_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3049_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3101__B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4515__326 vssd1 vssd1 vccd1 vccd1 _4515__326/HI net326 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4602__376 vssd1 vssd1 vccd1 vccd1 _4602__376/HI net376 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4676__444 vssd1 vssd1 vccd1 vccd1 _4676__444/HI net444 sky130_fd_sc_hd__conb_1
XFILLER_0_29_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2420_ net204 _0942_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4717__485 vssd1 vssd1 vccd1 vccd1 _4717__485/HI net485 sky130_fd_sc_hd__conb_1
XFILLER_0_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2351_ _1094_ _1097_ team_10_WB.instance_to_wrap.host_col\[2\] _0869_ vssd1 vssd1
+ vccd1 vccd1 _1127_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_62_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2282_ _0990_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4021_ clknet_leaf_49_wb_clk_i net583 _0068_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3485__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3805_ net278 vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
X_4785_ net182 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1997_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] net148 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1 vccd1 vccd1 _0752_
+ sky130_fd_sc_hd__o22a_1
X_3736_ net279 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout123_A _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3667_ net254 vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3872__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2618_ _1294_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] _1074_ vssd1 vssd1
+ vccd1 vccd1 _0006_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3598_ net287 vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2549_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\]
+ _1240_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\] vssd1 vssd1
+ vccd1 vccd1 _1241_ sky130_fd_sc_hd__o31a_2
XFILLER_0_122_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4219_ clknet_leaf_49_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[81\]
+ _0208_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[81\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3476__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3164__C1 _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
Xfanout291 net296 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_4
XFILLER_0_89_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1920_ net299 net2 vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4570_ net541 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3521_ net230 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2800__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3452_ team_10_WB.instance_to_wrap.host_row1\[54\] _1699_ net178 team_10_WB.instance_to_wrap.host_row2\[62\]
+ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2403_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ team_10_WB.instance_to_wrap.clock_div.count\[25\] team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__or4_1
XANTENNA__1924__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3383_ net302 _1758_ _1759_ net167 _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2334_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\] _0868_ vssd1 vssd1
+ vccd1 vccd1 _1110_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2265_ _1035_ _1040_ _1046_ _0949_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3458__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1940__A team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4004_ clknet_leaf_38_wb_clk_i _0492_ net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2130__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2196_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _0801_ _0978_ _0979_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout240_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4768_ net181 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3719_ net254 vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
X_4699_ net467 vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
XFILLER_0_120_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2011__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold11 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold22 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\] vssd1 vssd1 vccd1 vccd1
+ net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\] vssd1 vssd1 vccd1
+ vccd1 net585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 team_10_WB.instance_to_wrap.host_row1\[43\] vssd1 vssd1 vccd1 vccd1 net596
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3449__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 team_10_WB.instance_to_wrap.host_row1\[64\] vssd1 vssd1 vccd1 vccd1 net607
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_10_WB.instance_to_wrap.message_reg.msg\[1\] vssd1 vssd1 vccd1 vccd1 net618
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _0615_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 team_10_WB.instance_to_wrap.host_row1\[66\] vssd1 vssd1 vccd1 vccd1 net640
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold99 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] vssd1 vssd1 vccd1
+ vccd1 net651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2975__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2050_ team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] net114 net138 net812 vssd1
+ vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3687__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2415__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2952_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] net161 _1478_ net210 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[4\] sky130_fd_sc_hd__o22a_1
XFILLER_0_2_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4608__382 vssd1 vssd1 vccd1 vccd1 _4608__382/HI net382 sky130_fd_sc_hd__conb_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1903_ team_10_WB.instance_to_wrap.uart_receiver.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _0827_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2883_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] _1465_ vssd1 vssd1 vccd1
+ vccd1 _1466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4622_ team_10_WB.instance_to_wrap.uart_transmitter.tx_serial vssd1 vssd1 vccd1 vccd1
+ net75 sky130_fd_sc_hd__buf_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4553_ net364 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3504_ net236 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
XANTENNA__3391__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4484_ clknet_leaf_49_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[41\]
+ _0467_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\]
+ sky130_fd_sc_hd__dfstp_1
X_4732__500 vssd1 vssd1 vccd1 vccd1 _4732__500/HI net500 sky130_fd_sc_hd__conb_1
X_3435_ team_10_WB.instance_to_wrap.host_row2\[69\] team_10_WB.instance_to_wrap.dispFSM.guesses\[45\]
+ net300 vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3366_ net207 _0817_ _1690_ _1403_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2317_ net226 _0848_ net194 team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1
+ vccd1 vccd1 _1093_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout190_A _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3297_ net637 _1677_ _1678_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout288_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2248_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] _0801_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2179_ team_10_WB.instance_to_wrap.correct\[0\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2006__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3373__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3220_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ _1630_ vssd1
+ vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3151_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] _1551_ _1579_ _1580_ vssd1 vssd1
+ vccd1 vccd1 _0497_ sky130_fd_sc_hd__o22a_1
X_2102_ team_10_WB.instance_to_wrap.dispFSM.guesses\[10\] net110 net134 net821 vssd1
+ vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__o22a_1
X_3082_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _1535_ net201 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[77\] sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2033_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] net141 net108 net755 vssd1 vssd1
+ vccd1 vccd1 _0746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3984_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[21\]
+ _0052_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2939__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2935_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] net149 net120 net792 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[40\] sky130_fd_sc_hd__o22a_1
XFILLER_0_134_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2866_ net845 _1454_ net174 vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4605_ net379 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2797_ team_10_WB.instance_to_wrap.lcdPlayer.currentState\[3\] net175 vssd1 vssd1
+ vccd1 vccd1 _1406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 team_10_WB.instance_to_wrap.clock_div.count\[18\] vssd1 vssd1 vccd1 vccd1
+ net852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1
+ net863 sky130_fd_sc_hd__dlygate4sd3_1
X_4536_ net347 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 team_10_WB.instance_to_wrap.gamelogic.setWord\[32\] vssd1 vssd1 vccd1 vccd1
+ net874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4467_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[24\]
+ _0450_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3418_ _1790_ _1793_ net301 vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4398_ clknet_leaf_0_wb_clk_i _0783_ _0381_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[35\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_input8_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ _1680_ _1718_ net177 _1728_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_119_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2943__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3355__A2 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2563__B1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2720_ team_10_WB.instance_to_wrap.clock_div.count\[7\] _1351_ vssd1 vssd1 vccd1
+ vccd1 _1353_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2651_ _1310_ _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2582_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] _1259_ _0901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4321_ clknet_leaf_12_wb_clk_i _0711_ _0310_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[44\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4252_ clknet_leaf_52_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[8\]
+ _0241_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout109 net111 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3203_ _1619_ _1611_ _1618_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__and3b_1
X_4183_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[45\]
+ _0172_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[45\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3134_ _1563_ _1564_ net218 _0906_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_39_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3065_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2016_ net4 _0887_ _0892_ net225 vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__or4b_2
XFILLER_0_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3967_ clknet_leaf_42_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[4\]
+ _0035_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2918_ net676 net154 net124 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[23\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3898_ net262 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2849_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\] _1442_ vssd1 vssd1
+ vccd1 vccd1 _1445_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold130 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold141 team_10_WB.instance_to_wrap.dispFSM.guesses\[15\] vssd1 vssd1 vccd1 vccd1
+ net693 sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ net330 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xhold152 _0698_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 team_10_WB.instance_to_wrap.clock_div.count\[24\] vssd1 vssd1 vccd1 vccd1
+ net715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold174 team_10_WB.instance_to_wrap.host_row1\[49\] vssd1 vssd1 vccd1 vccd1 net726
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold185 team_10_WB.instance_to_wrap.clock_div.count\[3\] vssd1 vssd1 vccd1 vccd1
+ net737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold196 _0738_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4628__396 vssd1 vssd1 vccd1 vccd1 _4628__396/HI net396 sky130_fd_sc_hd__conb_1
XFILLER_0_77_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3009__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3821_ net250 vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3695__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3752_ net280 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2703_ net222 net218 net299 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__mux2_1
XFILLER_0_43_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3683_ net295 vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2634_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ _1083_ _1075_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__o31a_1
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2565_ _0974_ _1251_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4304_ clknet_leaf_15_wb_clk_i _0694_ _0293_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2496_ net224 _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4235_ clknet_leaf_31_wb_clk_i _0648_ _0224_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4166_ clknet_leaf_40_wb_clk_i _0635_ _0155_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3117_ net701 net5 _1548_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__mux2_1
X_4097_ clknet_leaf_8_wb_clk_i _0568_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout270_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3048_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _1518_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[60\] sky130_fd_sc_hd__mux2_1
XANTENNA__3170__A_N _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4554__365 vssd1 vssd1 vccd1 vccd1 _4554__365/HI net365 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2350_ _1124_ _1125_ _1099_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2281_ _1012_ _1061_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4020_ clknet_leaf_50_wb_clk_i net581 _0067_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2460__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3804_ net292 vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4784_ net181 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
X_1996_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _0874_ _0884_ net156 vssd1
+ vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3735_ net279 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__inv_2
X_4497__308 vssd1 vssd1 vccd1 vccd1 _4497__308/HI net308 sky130_fd_sc_hd__conb_1
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3666_ net271 vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout116_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2617_ _0830_ _1116_ _1119_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4538__349 vssd1 vssd1 vccd1 vccd1 _4538__349/HI net349 sky130_fd_sc_hd__conb_1
XFILLER_0_11_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3597_ net272 vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2548_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2920__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2479_ net614 net131 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4218_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[80\]
+ _0207_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[80\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4149_ clknet_leaf_9_wb_clk_i _0620_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2009__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4699__467 vssd1 vssd1 vccd1 vccd1 _4699__467/HI net467 sky130_fd_sc_hd__conb_1
XFILLER_0_19_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2911__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3467__A1 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout270 net274 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_4
Xfanout281 net297 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_2
Xfanout292 net296 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_4
XFILLER_0_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4643__411 vssd1 vssd1 vccd1 vccd1 _4643__411/HI net411 sky130_fd_sc_hd__conb_1
XFILLER_0_130_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3520_ net230 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3451_ net69 net175 _1825_ net227 vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2402_ team_10_WB.instance_to_wrap.clock_div.count\[27\] team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ team_10_WB.instance_to_wrap.clock_div.count\[29\] team_10_WB.instance_to_wrap.clock_div.count\[28\]
+ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__or4_1
XFILLER_0_81_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3382_ net206 _1690_ _1752_ net229 _1403_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2333_ _0810_ _0843_ _0855_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2264_ _1038_ _1039_ _1041_ _1043_ _1045_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4003_ clknet_leaf_38_wb_clk_i _0491_ net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2195_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _0802_ _0981_ _0983_ vssd1
+ vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2433__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout233_A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4767_ net181 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
X_1979_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3718_ net257 vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4698_ net466 vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
XFILLER_0_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3649_ net264 vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2011__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_10_WB.instance_to_wrap.host_row1\[61\] vssd1 vssd1 vccd1 vccd1 net564
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[5\] vssd1 vssd1 vccd1
+ vccd1 net575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold34 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[1\] vssd1 vssd1
+ vccd1 vccd1 net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 team_10_WB.instance_to_wrap.host_row1\[70\] vssd1 vssd1 vccd1 vccd1 net597
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_10_WB.instance_to_wrap.host_row1\[76\] vssd1 vssd1 vccd1 vccd1 net608
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_10_WB.instance_to_wrap.message_reg.msg\[7\] vssd1 vssd1 vccd1 vccd1 net619
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 team_10_WB.instance_to_wrap.host_row1\[67\] vssd1 vssd1 vccd1 vccd1 net630
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold89 team_10_WB.instance_to_wrap.host_row1\[50\] vssd1 vssd1 vccd1 vccd1 net641
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3385__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_9 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2951_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] net160 _1478_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[3\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_1902_ net199 vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2882_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] net221 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4621_ net392 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_72_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3376__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552_ net363 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_108_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3503_ net236 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4483_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[40\]
+ _0466_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_29_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3434_ team_10_WB.instance_to_wrap.host_row2\[85\] team_10_WB.instance_to_wrap.dispFSM.guesses\[61\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3365_ team_10_WB.instance_to_wrap.host_row2\[65\] team_10_WB.instance_to_wrap.dispFSM.guesses\[41\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2316_ net222 net223 _0850_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__and3b_1
X_3296_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ _1674_ net295 vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _0793_ net209 _0802_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] _1028_
+ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout183_A _0995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2178_ _0968_ team_10_WB.instance_to_wrap.correct\[1\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3118__A team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_124_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_102_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3358__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4755__523 vssd1 vssd1 vccd1 vccd1 _4755__523/HI net523 sky130_fd_sc_hd__conb_1
XFILLER_0_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3150_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] _1278_ _1568_ vssd1 vssd1 vccd1
+ vccd1 _1580_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2101_ team_10_WB.instance_to_wrap.dispFSM.guesses\[11\] net112 net140 net754 vssd1
+ vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__o22a_1
X_3081_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2032_ net193 _0903_ net136 vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3983_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[20\]
+ _0051_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2934_ net684 net154 net124 net729 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[39\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2865_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] _1454_ vssd1 vssd1
+ vccd1 vccd1 _1455_ sky130_fd_sc_hd__and2_1
XANTENNA__3349__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4604_ net378 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2796_ _1405_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4535_ net346 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_108_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold301 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] vssd1 vssd1 vccd1
+ vccd1 net853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] vssd1 vssd1 vccd1 vccd1
+ net864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold323 team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\] vssd1 vssd1 vccd1 vccd1
+ net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4466_ clknet_leaf_46_wb_clk_i net677 _0449_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3417_ team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] _1715_ _1791_ _1792_ vssd1
+ vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4397_ clknet_leaf_4_wb_clk_i _0782_ _0380_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3348_ team_10_WB.instance_to_wrap.host_row2\[64\] team_10_WB.instance_to_wrap.dispFSM.guesses\[40\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__mux2_1
X_3279_ net730 _1664_ net227 vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3401__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2017__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold310_A team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4739__507 vssd1 vssd1 vccd1 vccd1 _4739__507/HI net507 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4570__541 vssd1 vssd1 vccd1 vccd1 net541 _4570__541/LO sky130_fd_sc_hd__conb_1
XFILLER_0_25_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2251__B1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2650_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ _1224_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2581_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\] _0904_ _0906_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4320_ clknet_leaf_14_wb_clk_i _0710_ _0309_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[43\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_23_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4251_ clknet_leaf_52_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[7\]
+ _0240_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3202_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\]
+ _1392_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4182_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[44\]
+ _0171_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[44\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3133_ net216 _0905_ _1562_ _0907_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_78_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3064_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] _1526_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\] sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2015_ _0887_ _0892_ net225 vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3966_ clknet_leaf_44_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[3\]
+ _0034_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout146_A _0862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2917_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\] net151 net122 net828
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[22\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3897_ net259 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2848_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\] _1442_ vssd1 vssd1
+ vccd1 vccd1 _1444_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2779_ net863 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\] vssd1 vssd1 vccd1
+ vccd1 _1389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4202__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\] vssd1 vssd1 vccd1
+ vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ net329 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xhold131 team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs vssd1 vssd1 vccd1 vccd1 net683
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold142 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\] vssd1 vssd1 vccd1
+ vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold153 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\] vssd1 vssd1 vccd1 vccd1
+ net705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] vssd1 vssd1 vccd1 vccd1
+ net716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_10_WB.instance_to_wrap.dispFSM.guesses\[69\] vssd1 vssd1 vccd1 vccd1
+ net727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] vssd1 vssd1 vccd1 vccd1
+ net738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4449_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[6\]
+ _0432_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xhold197 team_10_WB.instance_to_wrap.dispFSM.guesses\[11\] vssd1 vssd1 vccd1 vccd1
+ net749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3131__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3820_ net259 vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__inv_2
XANTENNA__3016__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2224__A0 team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3751_ net279 vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2702_ net223 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] net299 vssd1
+ vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3682_ net249 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__inv_2
XANTENNA__1983__C1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2633_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] _1285_ _1290_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1300_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2564_ _1059_ _1250_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1
+ vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4303_ clknet_leaf_30_wb_clk_i _0693_ _0292_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\]
+ sky130_fd_sc_hd__dfstp_1
X_2495_ net229 _1177_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4234_ clknet_leaf_34_wb_clk_i _0647_ _0223_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4165_ clknet_leaf_40_wb_clk_i _0634_ _0154_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3116_ net666 net4 _1548_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4096_ clknet_leaf_8_wb_clk_i _0567_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3047_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout263_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4660__428 vssd1 vssd1 vccd1 vccd1 _4660__428/HI net428 sky130_fd_sc_hd__conb_1
XFILLER_0_33_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3949_ clknet_leaf_38_wb_clk_i _0012_ net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701__469 vssd1 vssd1 vccd1 vccd1 _4701__469/HI net469 sky130_fd_sc_hd__conb_1
XFILLER_0_89_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2280_ net215 _0952_ _1023_ _1060_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3803_ net272 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4783_ net182 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1995_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] net145 vssd1 vssd1
+ vccd1 vccd1 _0884_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3734_ net291 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1956__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3665_ net288 vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1971__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2616_ _0015_ _0012_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[2\]
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout109_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3596_ net269 vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3173__A1 _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2547_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _1239_ sky130_fd_sc_hd__and3b_1
XFILLER_0_80_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2478_ net592 net128 _1189_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__o22a_1
X_4217_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[79\]
+ _0206_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[79\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3476__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ clknet_leaf_9_wb_clk_i _0619_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_97_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4079_ clknet_leaf_36_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[10\]
+ _0099_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2987__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2025__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4521__332 vssd1 vssd1 vccd1 vccd1 _4521__332/HI net332 sky130_fd_sc_hd__conb_1
XFILLER_0_110_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1864__A team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3164__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input39_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 net265 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_4
Xfanout271 net273 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_4
Xfanout282 net286 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout293 net295 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4682__450 vssd1 vssd1 vccd1 vccd1 _4682__450/HI net450 sky130_fd_sc_hd__conb_1
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2978__B2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4723__491 vssd1 vssd1 vccd1 vccd1 _4723__491/HI net491 sky130_fd_sc_hd__conb_1
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3465__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3450_ _1781_ _1820_ _1824_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2401_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ _1160_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or4_1
X_3381_ team_10_WB.instance_to_wrap.host_row1\[58\] team_10_WB.instance_to_wrap.dispFSM.msg\[2\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2332_ _0843_ net194 _0810_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2263_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0800_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ _0790_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3458__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4002_ clknet_leaf_41_wb_clk_i _0490_ net244 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2194_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _0801_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ _0795_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2969__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4505__316 vssd1 vssd1 vccd1 vccd1 _4505__316/HI net316 sky130_fd_sc_hd__conb_1
XFILLER_0_16_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4766_ net180 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1978_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3717_ net252 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4697_ net465 vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
XFILLER_0_31_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3648_ net269 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3579_ net269 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold13 team_10_WB.instance_to_wrap.message_reg.msg\[5\] vssd1 vssd1 vccd1 vccd1 net565
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1
+ net576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\] vssd1 vssd1 vccd1 vccd1
+ net587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_10_WB.instance_to_wrap.host_row1\[51\] vssd1 vssd1 vccd1 vccd1 net598
+ sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_10_WB.instance_to_wrap.host_row1\[71\] vssd1 vssd1 vccd1 vccd1 net609
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _0526_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold79 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] vssd1 vssd1 vccd1
+ vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4666__434 vssd1 vssd1 vccd1 vccd1 _4666__434/HI net434 sky130_fd_sc_hd__conb_1
XFILLER_0_97_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3082__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4707__475 vssd1 vssd1 vccd1 vccd1 _4707__475/HI net475 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2896__B1 _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2950_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\] net161 _1478_ net212 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[2\] sky130_fd_sc_hd__o22a_1
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _0825_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2881_ _1222_ _1464_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_70_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4620_ net391 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_115_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4551_ net362 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3502_ net236 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4482_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[39\]
+ _0465_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3433_ team_10_WB.instance_to_wrap.host_row1\[69\] net301 _1703_ vssd1 vssd1 vccd1
+ vccd1 _1808_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3364_ _1738_ _1742_ _1736_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2315_ _0868_ _1090_ net4 vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__or3b_1
X_3295_ net295 _1676_ _1677_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _0804_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_75_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2177_ _0936_ _0962_ _0967_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3367__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4749_ net517 vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__buf_2
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_12_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2973__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2030__A1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2869__B1 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2100_ team_10_WB.instance_to_wrap.dispFSM.guesses\[12\] net115 net138 net854 vssd1
+ vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__o22a_1
X_3080_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] _1534_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[76\] sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2031_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _0886_ _0910_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__or4_2
XFILLER_0_136_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3982_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[19\]
+ _0050_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2933_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] net151 net122 net787
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[38\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2864_ _1454_ net174 _1453_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4603_ net377 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_32_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2795_ net228 _1404_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__nand2_2
XFILLER_0_25_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4621__392 vssd1 vssd1 vccd1 vccd1 _4621__392/HI net392 sky130_fd_sc_hd__conb_1
X_4534_ net345 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_48_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold302 team_10_WB.instance_to_wrap.dispFSM.guesses\[20\] vssd1 vssd1 vccd1 vccd1
+ net854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1
+ net865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] vssd1 vssd1 vccd1 vccd1
+ net876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4465_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[22\]
+ _0448_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_44_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1962__A team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3416_ team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] net169 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[12\]
+ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4396_ clknet_leaf_22_wb_clk_i _0781_ _0379_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3347_ _1682_ _1686_ _1688_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout293_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3278_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\]
+ _1663_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2229_ net768 net142 _0807_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3401__B net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2017__B net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input21_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3028__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2251__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2251__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2580_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\] _0906_ _1262_ _1263_
+ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4250_ clknet_leaf_52_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[6\]
+ _0239_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3201_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\]
+ _1391_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1
+ _1618_ sky130_fd_sc_hd__a31o_1
X_4181_ clknet_leaf_16_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\]
+ _0170_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[43\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3132_ _0890_ _0899_ _1259_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3063_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2014_ net2 net3 net4 net5 net300 vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__o41a_1
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3965_ clknet_leaf_44_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[2\]
+ _0033_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2916_ net657 net154 net124 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[21\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3896_ net263 vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout139_A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2847_ _1442_ _1443_ net174 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_33_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2778_ net557 _1388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[29\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold110 team_10_WB.instance_to_wrap.host_row1\[42\] vssd1 vssd1 vccd1 vccd1 net662
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold121 team_10_WB.instance_to_wrap.dispFSM.guesses\[45\] vssd1 vssd1 vccd1 vccd1
+ net673 sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ net328 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_41_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold132 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[47\] vssd1 vssd1 vccd1
+ vccd1 net684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[13\] vssd1 vssd1
+ vccd1 vccd1 net695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 team_10_WB.instance_to_wrap.host_row1\[46\] vssd1 vssd1 vccd1 vccd1 net706
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold165 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\] vssd1 vssd1 vccd1
+ vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold176 _0736_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ clknet_leaf_26_wb_clk_i net575 _0431_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold187 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold198 team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] vssd1 vssd1 vccd1 vccd1
+ net750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4379_ clknet_leaf_23_wb_clk_i _0764_ _0362_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2970__B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3998__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3249__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3750_ net291 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2701_ team_10_WB.instance_to_wrap.host_col\[0\] net220 net299 vssd1 vssd1 vccd1
+ vccd1 net78 sky130_fd_sc_hd__mux2_1
XFILLER_0_54_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3681_ net288 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2632_ net193 _1281_ _1298_ _0903_ _1299_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2563_ net751 _0948_ net133 vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4302_ clknet_leaf_30_wb_clk_i _0692_ _0291_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_107_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2494_ net632 net129 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] vssd1
+ vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__a22o_1
X_4233_ clknet_leaf_51_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[2\]
+ _0222_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4164_ clknet_leaf_44_wb_clk_i _0633_ _0153_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3115_ net671 net3 _1548_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4095_ clknet_leaf_9_wb_clk_i _0566_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3046_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _1517_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[59\] sky130_fd_sc_hd__mux2_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2463__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2463__B2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3948_ clknet_leaf_34_wb_clk_i _0011_ net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_50_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3412__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3879_ net283 vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3802_ net290 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4782_ net181 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1994_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] net146 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1 vccd1 _0754_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_111_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3733_ net239 vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3664_ net271 vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2615_ _1270_ _1282_ _1293_ _1275_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3595_ net269 vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2131__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2546_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2477_ net621 net131 _1185_ _1212_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4216_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[78\]
+ _0205_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[78\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4147_ clknet_leaf_12_wb_clk_i _0618_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4078_ clknet_leaf_36_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[9\]
+ _0098_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3029_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560__371 vssd1 vssd1 vccd1 vccd1 _4560__371/HI net371 sky130_fd_sc_hd__conb_1
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1880__A team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout250 net251 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_4
XANTENNA__2124__A0 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout261 net265 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_4
Xfanout283 net286 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_4
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4030__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2400_ team_10_WB.instance_to_wrap.clock_div.count\[11\] _1161_ _1162_ team_10_WB.instance_to_wrap.clock_div.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3380_ _1754_ _1755_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2331_ _0844_ net194 _0809_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__a21o_1
XANTENNA__3481__S net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2262_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] net212 vssd1 vssd1 vccd1
+ vccd1 _1044_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4001_ clknet_leaf_41_wb_clk_i _0489_ net244 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2193_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] _0804_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2969__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4544__355 vssd1 vssd1 vccd1 vccd1 _4544__355/HI net355 sky130_fd_sc_hd__conb_1
XFILLER_0_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4765_ net527 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_117_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1965__A team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1977_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] net147 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3716_ net252 vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout121_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4696_ net464 vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3647_ net258 vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3578_ net288 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2529_ net566 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0512_ sky130_fd_sc_hd__mux2_1
Xhold14 team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] vssd1 vssd1 vccd1 vccd1 net566
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold25 team_10_WB.instance_to_wrap.dispFSM.guesses\[7\] vssd1 vssd1 vccd1 vccd1 net577
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked vssd1 vssd1 vccd1 vccd1
+ net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_10_WB.instance_to_wrap.host_row1\[55\] vssd1 vssd1 vccd1 vccd1 net599
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] vssd1 vssd1 vccd1 vccd1 net610
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_10_WB.instance_to_wrap.host_row1\[54\] vssd1 vssd1 vccd1 vccd1 net621
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1875__A team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3385__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4528__339 vssd1 vssd1 vccd1 vccd1 _4528__339/HI net339 sky130_fd_sc_hd__conb_1
XFILLER_0_69_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1900_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] vssd1 vssd1 vccd1 vccd1
+ _0824_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2880_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] net1 _1463_ vssd1 vssd1 vccd1
+ vccd1 _1464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3376__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4550_ net361 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_108_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3501_ net237 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4481_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[38\]
+ _0464_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3432_ team_10_WB.instance_to_wrap.host_row1\[101\] net301 _1776_ _1806_ vssd1 vssd1
+ vccd1 vccd1 _1807_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_3363_ _1739_ _1740_ _1741_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__or3_1
XFILLER_0_110_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2314_ net222 net223 _0850_ _0818_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__o211ai_1
X_3294_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\]
+ _1672_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4689__457 vssd1 vssd1 vccd1 vccd1 _4689__457/HI net457 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _0800_ _0802_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__o221a_1
X_2176_ _0959_ _0960_ _0961_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4748_ net516 vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__buf_2
XFILLER_0_47_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4679_ net447 vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_2
XFILLER_0_120_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_4633__401 vssd1 vssd1 vccd1 vccd1 _4633__401/HI net401 sky130_fd_sc_hd__conb_1
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2973__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3358__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2566__B1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2030__A2 _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2030_ net193 _0903_ net141 vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3981_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[18\]
+ _0049_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2932_ net680 net155 _1472_ net672 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[37\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2863_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\]
+ _1450_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602_ net376 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_116_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2794_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[5\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4533_ net344 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
Xhold303 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold314 team_10_WB.instance_to_wrap.clock_div.count\[21\] vssd1 vssd1 vccd1 vccd1
+ net866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ net877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ clknet_leaf_32_wb_clk_i net658 _0447_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2309__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3415_ team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] _1701_ net166 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\]
+ _1771_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4395_ clknet_leaf_21_wb_clk_i _0780_ _0378_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3346_ _1722_ _1725_ _1713_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3277_ net626 _1661_ _1665_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout286_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2228_ net601 _1011_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2159_ _0924_ _0945_ _0951_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3401__C net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2984__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input14_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2251__A2 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output82_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3200_ _1612_ _1617_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4180_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[42\]
+ _0169_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[42\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3131_ net218 _1259_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__nor2_1
XANTENNA__2894__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3062_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] _1525_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[67\] sky130_fd_sc_hd__mux2_1
X_2013_ net300 net5 vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2490__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3964_ clknet_leaf_44_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[1\]
+ _0032_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2915_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\] net150 net121 net757
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[20\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3895_ net247 vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2846_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2777_ net732 _1388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[28\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold100 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[1\] vssd1 vssd1
+ vccd1 vccd1 net652 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4516_ net327 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
Xhold111 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout201_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 _0712_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 team_10_WB.instance_to_wrap.dispFSM.guesses\[37\] vssd1 vssd1 vccd1 vccd1
+ net685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold144 team_10_WB.instance_to_wrap.dispFSM.guesses\[21\] vssd1 vssd1 vccd1 vccd1
+ net696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2950__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 _0582_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4447_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[4\]
+ _0430_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\]
+ sky130_fd_sc_hd__dfstp_1
Xhold166 team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] vssd1 vssd1 vccd1 vccd1
+ net718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\] vssd1 vssd1 vccd1
+ vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold188 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1 net740
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold199 team_10_WB.instance_to_wrap.gamelogic.state\[0\] vssd1 vssd1 vccd1 vccd1
+ net751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4378_ clknet_leaf_25_wb_clk_i _0763_ _0361_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input6_A gpio_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3329_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _1682_ _1688_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4745__513 vssd1 vssd1 vccd1 vccd1 _4745__513/HI net513 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2466__C1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2233__A2 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2941__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3421__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3421__B2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2700_ _1342_ _1344_ _1238_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.tx_serial
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3680_ net272 vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2631_ _0911_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2562_ _0919_ _0972_ _1249_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4301_ clknet_leaf_13_wb_clk_i _0691_ _0290_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2493_ net636 net129 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] vssd1
+ vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4232_ clknet_leaf_51_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[1\]
+ _0221_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4163_ clknet_leaf_41_wb_clk_i _0632_ _0152_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3114_ net664 net2 _1548_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__mux2_1
X_4094_ clknet_leaf_9_wb_clk_i _0565_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2129__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3045_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2463__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout151_A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout249_A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3947_ clknet_leaf_21_wb_clk_i _0479_ _0021_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3878_ net283 vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1974__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1974__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2829_ _1411_ _1418_ _1426_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2923__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2439__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1878__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2914__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2221__B _1002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3801_ net281 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ net532 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1993_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] _0874_ _0883_ net156 vssd1
+ vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3732_ net240 vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1956__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3663_ net288 vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2614_ _0824_ _1287_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3594_ net284 vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2905__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2545_ net224 net553 _1216_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2381__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2476_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] net184 vssd1 vssd1 vccd1
+ vccd1 _1212_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4215_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[77\]
+ _0204_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[77\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout199_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4146_ clknet_leaf_8_wb_clk_i _0617_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4077_ clknet_leaf_35_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[8\]
+ _0097_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4781__532 vssd1 vssd1 vccd1 vccd1 _4781__532/HI net532 sky130_fd_sc_hd__conb_1
X_3028_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] _1508_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[50\] sky130_fd_sc_hd__mux2_1
XFILLER_0_78_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2009__D net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold209_A team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout240 net243 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_2
Xfanout251 net266 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_2
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout284 net286 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_4
Xfanout295 net296 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2216__B net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3388__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2060__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] _0819_ _0849_ vssd1
+ vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4650__418 vssd1 vssd1 vccd1 vccd1 _4650__418/HI net418 sky130_fd_sc_hd__conb_1
XFILLER_0_104_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2261_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] _0799_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\]
+ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3312__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4000_ clknet_leaf_41_wb_clk_i net644 net244 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2192_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _0802_ _0804_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4765__527 vssd1 vssd1 vccd1 vccd1 _4765__527/HI net527 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3379__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4622__A team_10_WB.instance_to_wrap.uart_transmitter.tx_serial vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4764_ net180 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1976_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _0874_ _0880_ net156 vssd1
+ vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3715_ net252 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4695_ net463 vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
XFILLER_0_16_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3646_ net261 vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3577_ net272 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2528_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold15 _0512_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] net195 _1185_
+ _1202_ net130 vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 _0674_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_10_WB.instance_to_wrap.message_reg.msg\[0\] vssd1 vssd1 vccd1 vccd1 net589
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold48 _0591_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 _0509_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4129_ clknet_leaf_28_wb_clk_i _0600_ _0128_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3701__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold326_A team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2896__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3500_ net235 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4480_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[37\]
+ _0463_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3431_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1805_ _1686_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3362_ team_10_WB.instance_to_wrap.host_row2\[49\] net168 _1708_ team_10_WB.instance_to_wrap.host_row1\[73\]
+ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__a22o_1
X_2313_ net226 _0848_ _0855_ net222 vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__o211a_1
X_3293_ net846 _1674_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2244_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0798_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4511__322 vssd1 vssd1 vccd1 vccd1 _4511__322/HI net322 sky130_fd_sc_hd__conb_1
XFILLER_0_75_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2175_ _0966_ team_10_WB.instance_to_wrap.correct\[2\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2137__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4747_ net515 vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__buf_2
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] net147 net119 net876 vssd1
+ vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4678_ net446 vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_2
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3629_ net247 vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4672__440 vssd1 vssd1 vccd1 vccd1 _4672__440/HI net440 sky130_fd_sc_hd__conb_1
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_99_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4713__481 vssd1 vssd1 vccd1 vccd1 _4713__481/HI net481 sky130_fd_sc_hd__conb_1
XFILLER_0_118_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2263__B1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3460__C1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2213__C net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2869__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3980_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[17\]
+ _0048_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2931_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] net150 net121 net762
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[36\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3451__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2862_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ _1448_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\] vssd1 vssd1 vccd1
+ vccd1 _1453_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4601_ net375 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_13_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2793_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] _1393_ _1395_ _1402_
+ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__or4_4
XFILLER_0_115_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4532_ net343 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_108_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4656__424 vssd1 vssd1 vccd1 vccd1 _4656__424/HI net424 sky130_fd_sc_hd__conb_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold304 team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1 vccd1 vccd1
+ net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold315 team_10_WB.instance_to_wrap.dispFSM.guesses\[41\] vssd1 vssd1 vccd1 vccd1
+ net867 sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[20\]
+ _0446_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_29_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 net878
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2309__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3414_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1704_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[68\]
+ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4394_ clknet_leaf_47_wb_clk_i _0779_ _0377_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4043__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3345_ _1716_ _1723_ _1724_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3276_ net294 _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2227_ team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] _1009_ _1010_ _0808_
+ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout181_A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2493__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2158_ net215 net214 _0947_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2089_ team_10_WB.instance_to_wrap.dispFSM.guesses\[31\] net143 net108 net687 vssd1
+ vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2984__B _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2236__B1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3130_ _1286_ _1554_ _1560_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3061_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2012_ net300 net5 vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__and2_1
XANTENNA__2475__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3963_ clknet_leaf_44_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[0\]
+ _0031_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2914_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\] net150 net121 net770
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[19\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3894_ net248 vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1986__C1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2845_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1442_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2776_ team_10_WB.instance_to_wrap.clock_div.count\[27\] team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ team_10_WB.instance_to_wrap.clock_div.count\[28\] _1384_ vssd1 vssd1 vccd1 vccd1
+ _1388_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4515_ net326 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
Xhold101 team_10_WB.instance_to_wrap.host_row1\[68\] vssd1 vssd1 vccd1 vccd1 net653
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 net664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold123 team_10_WB.instance_to_wrap.clock_div.count\[4\] vssd1 vssd1 vccd1 vccd1
+ net675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 team_10_WB.instance_to_wrap.host_row1\[69\] vssd1 vssd1 vccd1 vccd1 net686
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold145 _0688_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2150__A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold156 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\] vssd1 vssd1 vccd1
+ vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2950__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4446_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[3\]
+ _0429_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\]
+ sky130_fd_sc_hd__dfstp_1
Xhold167 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\] vssd1 vssd1 vccd1
+ vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4377_ clknet_leaf_3_wb_clk_i _0762_ _0360_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2702__A1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3328_ _1697_ _1707_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3259_ net293 _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2941__A1 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2630_ _0886_ _0909_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2561_ net215 net214 _0947_ _1034_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__a41o_1
XFILLER_0_45_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4300_ clknet_leaf_29_wb_clk_i net688 _0289_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2492_ net662 net132 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\] vssd1
+ vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4231_ clknet_leaf_51_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[0\]
+ _0220_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4162_ clknet_leaf_41_wb_clk_i _0631_ _0151_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3113_ net663 net216 _1548_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__mux2_1
X_4093_ clknet_leaf_9_wb_clk_i _0564_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3044_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] _1516_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[58\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2999__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout144_A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3946_ clknet_leaf_22_wb_clk_i _0478_ _0020_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3412__A2 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3877_ net249 vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2828_ _1409_ _0513_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2759_ team_10_WB.instance_to_wrap.clock_div.count\[21\] _1376_ vssd1 vssd1 vccd1
+ vccd1 _1378_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4429_ clknet_leaf_17_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[26\]
+ _0412_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3479__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3704__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2439__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3100__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3167__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2221__C _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3800_ net278 vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4780_ net182 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1992_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] net145 vssd1 vssd1
+ vccd1 vccd1 _0883_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3731_ net242 vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3662_ net258 vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2613_ _0016_ _0014_ _0015_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3593_ net269 vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2544_ team_10_WB.instance_to_wrap.host_col\[0\] _1237_ _1179_ vssd1 vssd1 vccd1
+ vccd1 _0484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2475_ net599 net129 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__a22o_1
X_4214_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[76\]
+ _0203_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[76\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4145_ clknet_leaf_16_wb_clk_i _0616_ _0144_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4076_ clknet_leaf_35_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[7\]
+ _0096_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3027_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout261_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3929_ net255 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1920__A_N net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout230 net233 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_4
Xfanout252 net255 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_4
Xfanout263 net265 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout274 net297 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_2
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_4
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4567__538 vssd1 vssd1 vccd1 vccd1 net538 _4567__538/LO sky130_fd_sc_hd__conb_1
XANTENNA__3085__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2232__B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2899__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2260_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0800_ vssd1 vssd1 vccd1
+ vccd1 _1042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2191_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] team_10_WB.instance_to_wrap.gamelogic.letter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__xor2_1
X_4730__498 vssd1 vssd1 vccd1 vccd1 _4730__498/HI net498 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3076__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4763_ net181 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1975_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] net145 vssd1 vssd1 vccd1
+ vccd1 _0880_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3714_ net252 vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__inv_2
X_4694_ net462 vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
XFILLER_0_71_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3645_ net262 vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3576_ net260 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2527_ team_10_WB.instance_to_wrap.uart_receiver.state\[0\] team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] vssd1 vssd1 vccd1 vccd1 _1233_
+ sky130_fd_sc_hd__or3b_4
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2458_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] net183 vssd1 vssd1 vccd1
+ vccd1 _1202_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] vssd1 vssd1 vccd1 vccd1 net568
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold27 team_10_WB.instance_to_wrap.message_reg.msg\[4\] vssd1 vssd1 vccd1 vccd1 net579
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 team_10_WB.instance_to_wrap.message_reg.msg\[2\] vssd1 vssd1 vccd1 vccd1 net590
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_10_WB.instance_to_wrap.message_reg.state\[1\] vssd1 vssd1 vccd1 vccd1
+ net601 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _0844_ net682 _1158_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4128_ clknet_leaf_24_wb_clk_i _0599_ _0127_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3067__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4059_ clknet_leaf_7_wb_clk_i _0544_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2599__A_N _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input37_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3103__S net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3430_ net206 _0817_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3361_ team_10_WB.instance_to_wrap.host_row1\[49\] _1699_ net167 team_10_WB.instance_to_wrap.host_row1\[57\]
+ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__a22o_1
X_2312_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3292_ net645 _1672_ _1675_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2243_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] _0805_ vssd1 vssd1 vccd1
+ vccd1 _1025_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550__361 vssd1 vssd1 vccd1 vccd1 _4550__361/HI net361 sky130_fd_sc_hd__conb_1
XFILLER_0_79_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2174_ _0964_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3049__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2272__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4746_ net514 vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__buf_2
XFILLER_0_133_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1958_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[35\]
+ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4677_ net445 vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1889_ net855 vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3628_ net245 vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3559_ net275 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3288__B1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3712__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2263__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3460__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_90 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2998__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2213__D net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4493__304 vssd1 vssd1 vccd1 vccd1 _4493__304/HI net304 sky130_fd_sc_hd__conb_1
XFILLER_0_105_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4534__345 vssd1 vssd1 vccd1 vccd1 _4534__345/HI net345 sky130_fd_sc_hd__conb_1
XFILLER_0_101_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3279__B1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2930_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] net150 net121 net796
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[35\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2861_ net633 _1450_ _1452_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4600_ net552 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_0_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2792_ _1396_ _1400_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4531_ net342 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4695__463 vssd1 vssd1 vccd1 vccd1 _4695__463/HI net463 sky130_fd_sc_hd__conb_1
XFILLER_0_124_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold305 team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1 vssd1 vccd1 vccd1
+ net857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold316 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\] vssd1 vssd1 vccd1
+ vccd1 net868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4462_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[19\]
+ _0445_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3413_ team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] net179 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4393_ clknet_leaf_4_wb_clk_i _0778_ _0376_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_106_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2420__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3344_ team_10_WB.instance_to_wrap.dispFSM.guesses\[0\] _1717_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[64\]
+ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3275_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] _1661_ vssd1 vssd1 vccd1
+ vccd1 _1664_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3532__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2226_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _1010_ sky130_fd_sc_hd__or3b_1
XFILLER_0_119_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2157_ net214 _0916_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2088_ team_10_WB.instance_to_wrap.dispFSM.guesses\[24\] net113 net137 net721 vssd1
+ vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2245__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4729_ net497 vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_2
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3707__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4518__329 vssd1 vssd1 vccd1 vccd1 _4518__329/HI net329 sky130_fd_sc_hd__conb_1
XFILLER_0_40_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1897__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3433__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4605__379 vssd1 vssd1 vccd1 vccd1 _4605__379/HI net379 sky130_fd_sc_hd__conb_1
X_4679__447 vssd1 vssd1 vccd1 vccd1 _4679__447/HI net447 sky130_fd_sc_hd__conb_1
XFILLER_0_129_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3617__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output68_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3060_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] _1524_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[66\] sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2011_ net300 net4 vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3962_ clknet_leaf_34_wb_clk_i _0482_ _0030_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3424__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2913_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\] net150 net121 net779
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[18\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3893_ net260 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2844_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] net585 _1441_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2775_ team_10_WB.instance_to_wrap.clock_div.count\[27\] _1386_ net731 vssd1 vssd1
+ vccd1 vccd1 _1387_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4514_ net325 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_108_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2431__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold102 team_10_WB.instance_to_wrap.host_row1\[74\] vssd1 vssd1 vccd1 vccd1 net654
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] vssd1 vssd1 vccd1 vccd1
+ net665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold124 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\] vssd1 vssd1 vccd1
+ vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold135 team_10_WB.instance_to_wrap.dispFSM.guesses\[23\] vssd1 vssd1 vccd1 vccd1
+ net687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4445_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[2\]
+ _0428_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 team_10_WB.instance_to_wrap.dispFSM.guesses\[13\] vssd1 vssd1 vccd1 vccd1
+ net698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 team_10_WB.instance_to_wrap.dispFSM.guesses\[5\] vssd1 vssd1 vccd1 vccd1
+ net709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[15\] vssd1 vssd1
+ vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold179 team_10_WB.instance_to_wrap.clock_div.count\[28\] vssd1 vssd1 vccd1 vccd1
+ net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4376_ clknet_leaf_46_wb_clk_i _0761_ _0359_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__3360__C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3327_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _0817_ vssd1 vssd1 vccd1
+ vccd1 _1707_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout291_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3258_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] _1651_ vssd1 vssd1 vccd1
+ vccd1 _1653_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2466__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2209_ net591 _0996_ _0992_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__o21a_1
X_3189_ net293 net176 _1610_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__or3_2
XFILLER_0_55_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3415__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1977__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2941__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3351__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1968__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4499__310 vssd1 vssd1 vccd1 vccd1 _4499__310/HI net310 sky130_fd_sc_hd__conb_1
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2955__A1_N _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2560_ _0973_ _1248_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2932__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2491_ net596 net132 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] vssd1
+ vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__a22o_1
X_4230_ clknet_leaf_57_wb_clk_i _0646_ _0219_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4161_ clknet_leaf_41_wb_clk_i _0630_ _0150_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3112_ net624 net217 _1548_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__mux2_1
X_4092_ clknet_leaf_9_wb_clk_i _0563_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3043_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2426__A _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3945_ clknet_leaf_0_wb_clk_i _0477_ _0019_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3876_ net260 vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2827_ _1407_ _1418_ _1429_ _1427_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2758_ net866 _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2923__A2 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2689_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] _1336_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_111_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4428_ clknet_leaf_16_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[25\]
+ _0411_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2136__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4359_ clknet_leaf_10_wb_clk_i _0002_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_5_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3720__A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2914__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1991_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3730_ net240 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3661_ net262 vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2612_ net193 _0909_ _1292_ _1290_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3592_ net284 vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__inv_2
X_4735__503 vssd1 vssd1 vccd1 vccd1 _4735__503/HI net503 sky130_fd_sc_hd__conb_1
XFILLER_0_109_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2905__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2543_ _0819_ team_10_WB.instance_to_wrap.host_col\[0\] _0851_ vssd1 vssd1 vccd1
+ vccd1 _1237_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2474_ net622 net128 _1211_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__o21a_1
X_4618__389 vssd1 vssd1 vccd1 vccd1 _4618__389/HI net389 sky130_fd_sc_hd__conb_1
X_4213_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[75\]
+ _0202_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[75\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4144_ clknet_leaf_24_wb_clk_i net629 _0143_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4075_ clknet_leaf_35_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[6\]
+ _0095_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3026_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _1507_ net199 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[49\] sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1995__A team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3397__A2 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3928_ net256 vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3859_ net283 vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3715__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2109__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout220 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\] vssd1 vssd1 vccd1
+ vccd1 net220 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_4
Xfanout253 net255 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_4
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout286 net297 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3388__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2060__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2190_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] net209 vssd1 vssd1 vccd1
+ vccd1 _0979_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3379__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4762_ net180 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1974_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] net147 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\]
+ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4624__393 vssd1 vssd1 vccd1 vccd1 _4624__393/HI net393 sky130_fd_sc_hd__conb_1
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3713_ net252 vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2423__B _1184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4693_ net461 vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_2
XFILLER_0_132_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3644_ net248 vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3575_ net285 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2526_ net589 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1
+ vccd1 vccd1 _0519_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2457_ net604 net128 _1201_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold17 _0507_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold28 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] vssd1 vssd1 vccd1 vccd1 net580
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 team_10_WB.instance_to_wrap.gamelogic.red vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ net5 net735 _1158_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4127_ clknet_leaf_15_wb_clk_i _0598_ _0126_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3270__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4058_ clknet_leaf_7_wb_clk_i _0543_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3009_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] net186 vssd1 vssd1 vccd1
+ vccd1 _1499_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3360_ team_10_WB.instance_to_wrap.host_row2\[57\] net178 net165 team_10_WB.instance_to_wrap.host_row2\[73\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2311_ _0841_ _1069_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__or3b_2
X_3291_ net295 _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2242_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2173_ _0959_ _0962_ _0963_ _0937_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2272__A2 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4745_ net513 vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__buf_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] net147 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4676_ net444 vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_2
XFILLER_0_31_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1888_ net216 vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3627_ net245 vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3265__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2416__A_N _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3558_ net275 vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__inv_2
X_2509_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] net221 _1225_ vssd1
+ vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3489_ net254 vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2263__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4640__408 vssd1 vssd1 vccd1 vccd1 _4640__408/HI net408 sky130_fd_sc_hd__conb_1
XFILLER_0_81_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_80 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_91 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2971__B1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3451__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2860_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] _1450_ net174
+ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2791_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4530_ net341 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4461_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[18\]
+ _0444_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold306 team_10_WB.instance_to_wrap.clock_div.count\[26\] vssd1 vssd1 vccd1 vccd1
+ net858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\] vssd1 vssd1 vccd1
+ vccd1 net869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3412_ team_10_WB.instance_to_wrap.host_row1\[60\] _1704_ _1708_ team_10_WB.instance_to_wrap.host_row1\[76\]
+ _1787_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4392_ clknet_leaf_47_wb_clk_i _0777_ _0375_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3343_ team_10_WB.instance_to_wrap.dispFSM.guesses\[24\] net168 net167 team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ net229 vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3274_ net638 _1660_ _1662_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2225_ _0808_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__or3b_1
XFILLER_0_20_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3024__S net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2156_ _0949_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2087_ team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] net109 net135 net837 vssd1
+ vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout167_A _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2245__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2989_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\] net160 _1491_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[27\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4728_ net496 vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4659_ net427 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_115_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4557__368 vssd1 vssd1 vccd1 vccd1 _4557__368/HI net368 sky130_fd_sc_hd__conb_1
XFILLER_0_102_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2236__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4501__312 vssd1 vssd1 vccd1 vccd1 _4501__312/HI net312 sky130_fd_sc_hd__conb_1
XFILLER_0_1_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold8_A team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2010_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\] net217 net219 net220
+ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ clknet_leaf_34_wb_clk_i _0481_ _0029_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_4662__430 vssd1 vssd1 vccd1 vccd1 _4662__430/HI net430 sky130_fd_sc_hd__conb_1
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2912_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\] net149 net120 net790
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[17\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3892_ net264 vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1986__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2843_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] net585 net174
+ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4703__471 vssd1 vssd1 vccd1 vccd1 _4703__471/HI net471 sky130_fd_sc_hd__conb_1
XFILLER_0_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2774_ net660 _1386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[27\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2935__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4513_ net324 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_79_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold114 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 net666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold125 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[23\] vssd1 vssd1
+ vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4444_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[1\]
+ _0427_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\]
+ sky130_fd_sc_hd__dfstp_1
Xhold136 _0690_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold147 team_10_WB.instance_to_wrap.dispFSM.guesses\[47\] vssd1 vssd1 vccd1 vccd1
+ net699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold158 team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\] vssd1 vssd1 vccd1 vccd1
+ net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\] vssd1 vssd1 vccd1 vccd1
+ net721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4375_ clknet_leaf_2_wb_clk_i _0760_ _0358_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3360__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3326_ team_10_WB.instance_to_wrap.host_row2\[80\] net171 net168 team_10_WB.instance_to_wrap.host_row2\[48\]
+ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3257_ _1651_ _1652_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2208_ _0946_ _0995_ _0990_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3188_ net293 net176 _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__nor3_4
XFILLER_0_69_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2466__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2139_ net133 _0934_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3718__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3103__A0 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2457__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4646__414 vssd1 vssd1 vccd1 vccd1 _4646__414/HI net414 sky130_fd_sc_hd__conb_1
XFILLER_0_19_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3406__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2917__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2490_ net615 net131 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] vssd1
+ vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3342__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4160_ clknet_leaf_42_wb_clk_i net649 _0149_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3111_ net647 net219 _1548_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__mux2_1
X_4091_ clknet_leaf_9_wb_clk_i _0562_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3042_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] _1515_ net199 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[57\] sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2448__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3944_ clknet_leaf_57_wb_clk_i _0476_ _0018_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1959__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3875_ net260 vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3538__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2826_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2757_ _1375_ _1376_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[20\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2688_ _1336_ _1337_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_1305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4427_ clknet_leaf_16_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[24\]
+ _0410_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ clknet_leaf_10_wb_clk_i _0001_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _0815_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1679_ vssd1 vssd1
+ vccd1 vccd1 _1690_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ clknet_leaf_12_wb_clk_i _0679_ _0278_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_119_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2439__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3100__A3 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2072__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3911__A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4150__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1990_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] net144 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3660_ net272 vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2611_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ _1291_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3591_ net285 vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2366__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2542_ net223 _1068_ _1179_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2473_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] net195 _1185_
+ _1210_ net130 vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590__549 vssd1 vssd1 vccd1 vccd1 net549 _4590__549/LO sky130_fd_sc_hd__conb_1
X_4212_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[74\]
+ _0201_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[74\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4143_ clknet_leaf_3_wb_clk_i _0614_ _0142_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4074_ clknet_leaf_36_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[5\]
+ _0094_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3025_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\]
+ net185 vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout247_A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3927_ net241 vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3858_ net282 vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2809_ net227 _1414_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3789_ net278 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout210 team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1
+ net210 sky130_fd_sc_hd__buf_4
Xfanout221 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\] vssd1 vssd1 vccd1
+ vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_4
Xfanout243 net266 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_4
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout276 net297 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_4
Xfanout287 net297 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_4
Xfanout298 net7 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2045__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2899__A2 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2520__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4761_ net526 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2036__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1973_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0874_ _0879_ net156 vssd1
+ vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3712_ net298 vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4692_ net460 vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3643_ net259 vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3574_ net287 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4046__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2525_ net618 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1
+ vccd1 vccd1 _0520_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3027__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2456_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] net195 team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\]
+ net126 net130 vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold18 team_10_WB.instance_to_wrap.message_reg.msg\[6\] vssd1 vssd1 vccd1 vccd1 net570
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold29 _0505_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0856_ vssd1 vssd1 vccd1
+ vccd1 _1158_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4126_ clknet_leaf_27_wb_clk_i _0597_ _0125_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4057_ clknet_leaf_6_wb_clk_i _0542_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3008_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\] net183 _1498_ net201
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[40\] sky130_fd_sc_hd__o211a_1
XFILLER_0_78_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3472__C1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3726__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4573__544 vssd1 vssd1 vccd1 vccd1 net544 _4573__544/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2310_ team_10_WB.instance_to_wrap.host_col\[0\] _0859_ _0864_ vssd1 vssd1 vccd1
+ vccd1 _1086_ sky130_fd_sc_hd__or3b_1
X_3290_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] _1668_ vssd1 vssd1 vccd1 vccd1
+ _1674_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2241_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] _1022_ _1013_ _1015_
+ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__or4b_2
XFILLER_0_40_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2172_ _0959_ _0962_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4744_ net512 vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__buf_2
X_1956_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0874_ _0876_ net158 vssd1
+ vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4675_ net443 vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_2
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1887_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 _0811_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3626_ net245 vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2980__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout112_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3557_ net275 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2508_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] _1224_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__o21a_2
X_3488_ net252 vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2439_ net654 net131 net125 team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4109_ clknet_leaf_18_wb_clk_i _0580_ _0108_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3460__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4720__488 vssd1 vssd1 vccd1 vccd1 _4720__488/HI net488 sky130_fd_sc_hd__conb_1
XANTENNA_70 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_81 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_92 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input42_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2487__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3436__C1 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3451__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2254__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2790_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2270__A team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4460_ clknet_leaf_47_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[17\]
+ _0443_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2962__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 team_10_WB.instance_to_wrap.clock_div.count\[22\] vssd1 vssd1 vccd1 vccd1
+ net859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold318 team_10_WB.instance_to_wrap.dispFSM.guesses\[43\] vssd1 vssd1 vccd1 vccd1
+ net870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3411_ team_10_WB.instance_to_wrap.host_row2\[52\] net168 _1784_ _1786_ vssd1 vssd1
+ vccd1 vccd1 _1787_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4391_ clknet_leaf_1_wb_clk_i _0776_ _0374_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3342_ team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] net172 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[8\]
+ _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3273_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ vssd1 vssd1 vccd1 vccd1
+ _1663_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2224_ team_10_WB.EN_VAL_REG net41 _1008_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2155_ _0935_ _0948_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2086_ team_10_WB.instance_to_wrap.dispFSM.guesses\[26\] net110 net134 net818 vssd1
+ vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3040__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2988_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\] net160 _1491_ net212
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[26\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4727_ net495 vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_2
X_1939_ team_10_WB.instance_to_wrap.host_message_reg.Cstate team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] _0861_ vssd1 vssd1 vccd1 vccd1
+ _0862_ sky130_fd_sc_hd__or4_2
XFILLER_0_86_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3276__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2953__A1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4658_ net426 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3609_ net284 vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4589_ net548 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2469__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4540__351 vssd1 vssd1 vccd1 vccd1 _4540__351/HI net351 sky130_fd_sc_hd__conb_1
XFILLER_0_50_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ clknet_leaf_34_wb_clk_i _0480_ _0028_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2911_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\] net149 net120 net777
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[16\]
+ sky130_fd_sc_hd__o22a_1
X_3891_ net260 vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2842_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] net174 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[0\] sky130_fd_sc_hd__and2b_1
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2773_ _1385_ _1386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[26\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2935__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4512_ net323 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_87_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\] vssd1 vssd1 vccd1
+ vccd1 net656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold126 team_10_WB.instance_to_wrap.host_row1\[48\] vssd1 vssd1 vccd1 vccd1 net678
+ sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[0\]
+ _0426_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold137 team_10_WB.instance_to_wrap.dispFSM.guesses\[61\] vssd1 vssd1 vccd1 vccd1
+ net689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold148 _0714_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold159 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\] vssd1 vssd1 vccd1
+ vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4374_ clknet_leaf_20_wb_clk_i _0759_ _0357_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3325_ team_10_WB.instance_to_wrap.host_row1\[64\] _1703_ net167 team_10_WB.instance_to_wrap.host_row1\[56\]
+ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3256_ _0813_ _1650_ net293 vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ net192 _0993_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__or2_2
XFILLER_0_20_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _0814_ _1607_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__or3b_4
XFILLER_0_119_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2871__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2138_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ _0926_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2069_ team_10_WB.instance_to_wrap.dispFSM.guesses\[43\] net111 net136 net823 vssd1
+ vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__o22a_1
XANTENNA__3415__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4524__335 vssd1 vssd1 vccd1 vccd1 _4524__335/HI net335 sky130_fd_sc_hd__conb_1
XFILLER_0_130_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3351__A1 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3103__A1 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4611__385 vssd1 vssd1 vccd1 vccd1 _4611__385/HI net385 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4685__453 vssd1 vssd1 vccd1 vccd1 _4685__453/HI net453 sky130_fd_sc_hd__conb_1
XFILLER_0_73_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4726__494 vssd1 vssd1 vccd1 vccd1 _4726__494/HI net494 sky130_fd_sc_hd__conb_1
XFILLER_0_131_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1968__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output73_A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3110_ net643 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\] _1548_ vssd1
+ vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__mux2_1
X_4090_ clknet_leaf_9_wb_clk_i _0561_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3041_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\]
+ net185 vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4508__319 vssd1 vssd1 vccd1 vccd1 _4508__319/HI net319 sky130_fd_sc_hd__conb_1
XFILLER_0_8_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3943_ net298 vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3874_ net260 vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2825_ net228 _1412_ _1417_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2756_ team_10_WB.instance_to_wrap.clock_div.count\[19\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ _1372_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2687_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] _1334_ _1319_ vssd1
+ vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3554__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4426_ clknet_leaf_24_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[23\]
+ _0409_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2315__C_N net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4357_ clknet_leaf_10_wb_clk_i _0000_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net207 _1686_ _1688_
+ _1685_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ clknet_leaf_15_wb_clk_i _0678_ _0277_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_4669__437 vssd1 vssd1 vccd1 vccd1 _4669__437/HI net437 sky130_fd_sc_hd__conb_1
X_3239_ _1642_ _1611_ _1641_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__and3b_1
XFILLER_0_55_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3729__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4583__546 vssd1 vssd1 vccd1 vccd1 net546 _4583__546/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2262__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2610_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3590_ net249 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2541_ net222 _1236_ _1179_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2472_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] net183 vssd1 vssd1 vccd1
+ vccd1 _1210_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3093__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4211_ clknet_leaf_49_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[73\]
+ _0200_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[73\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4142_ clknet_leaf_15_wb_clk_i _0613_ _0141_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4073_ clknet_leaf_36_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[4\]
+ _0093_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3024_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] _1506_ net199 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[48\] sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3094__A3 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout142_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3926_ net241 vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3857_ net282 vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2808_ net207 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[2\] _1403_ vssd1
+ vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3788_ net292 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2739_ _1363_ _1364_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4409_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[6\]
+ _0392_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_4
Xfanout211 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1
+ net211 sky130_fd_sc_hd__clkbuf_4
Xfanout222 team_10_WB.instance_to_wrap.host_col\[2\] vssd1 vssd1 vccd1 vccd1 net222
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout244 net246 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_4
Xfanout255 net266 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout266 net298 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_4
Xfanout288 net297 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
Xfanout299 net300 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2257__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4760_ net181 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2036__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1972_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] net144 vssd1 vssd1 vccd1
+ vccd1 _0879_ sky130_fd_sc_hd__or2_1
X_3711_ net231 vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4691_ net459 vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_2
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3642_ net249 vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3573_ net272 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2524_ net590 _1231_ _1232_ net878 vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2455_ net607 net129 _1185_ _1200_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold19 team_10_WB.instance_to_wrap.host_row1\[62\] vssd1 vssd1 vccd1 vccd1 net571
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] _1084_ _1156_
+ _1157_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__o22a_1
X_4125_ clknet_leaf_16_wb_clk_i _0596_ _0124_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3043__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4631__399 vssd1 vssd1 vccd1 vccd1 _4631__399/HI net399 sky130_fd_sc_hd__conb_1
X_4056_ clknet_leaf_6_wb_clk_i _0541_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3007_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] net187 vssd1 vssd1 vccd1
+ vccd1 _1498_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3909_ net250 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2240_ _1016_ _1017_ _1019_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__or4b_1
XFILLER_0_104_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2171_ team_10_WB.instance_to_wrap.correct\[2\] team_10_WB.instance_to_wrap.gamelogic.rights\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3454__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4743_ net511 vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_2
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1955_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] net144 vssd1 vssd1 vccd1
+ vccd1 _0876_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4674_ net442 vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1886_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 _0810_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2450__B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3625_ net247 vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3556_ net232 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2507_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] _1223_ vssd1 vssd1
+ vccd1 vccd1 _1224_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3487_ net254 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
X_2438_ net670 net131 _1191_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__a221o_1
X_2369_ _0871_ _1143_ _1087_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__a21oi_1
X_4108_ clknet_leaf_11_wb_clk_i _0579_ _0107_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4039_ clknet_leaf_33_wb_clk_i _0524_ _0080_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_60 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_93 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input35_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2239__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3436__B1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1998__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2270__B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1 vccd1
+ vccd1 net860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 team_10_WB.instance_to_wrap.dispFSM.guesses\[9\] vssd1 vssd1 vccd1 vccd1
+ net871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3410_ team_10_WB.instance_to_wrap.host_row1\[68\] _1703_ net178 team_10_WB.instance_to_wrap.host_row2\[60\]
+ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4390_ clknet_leaf_0_wb_clk_i _0775_ _0373_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3341_ team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] _1701_ net178 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\]
+ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3272_ net294 _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2223_ net42 net40 net43 _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2154_ _0822_ net214 _0948_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2085_ team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] net112 net140 net802 vssd1
+ vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2445__B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1989__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2987_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] net162 _1491_ net213
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[25\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4726_ net494 vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_2
XFILLER_0_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1938_ _0840_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2953__A2 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4657_ net425 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_16_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1869_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] vssd1 vssd1 vccd1 vccd1
+ _0794_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3608_ net285 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4588_ net547 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_29_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3539_ net239 vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4059__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2636__A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3930__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3409__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2880__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2910_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\] net154 net124 net719
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[15\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2632__A1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2632__B2 _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3890_ net261 vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2841_ _1010_ _1238_ _1241_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4777__530 vssd1 vssd1 vccd1 vccd1 _4777__530/HI net530 sky130_fd_sc_hd__conb_1
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2772_ team_10_WB.instance_to_wrap.clock_div.count\[25\] team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ team_10_WB.instance_to_wrap.clock_div.count\[26\] _1382_ vssd1 vssd1 vccd1 vccd1
+ _1386_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4511_ net322 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold105 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\] vssd1 vssd1 vccd1
+ vccd1 net657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 team_10_WB.instance_to_wrap.clock_div.count\[0\] vssd1 vssd1 vccd1 vccd1
+ net668 sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[39\]
+ _0425_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold138 _0728_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\] vssd1 vssd1 vccd1
+ vccd1 net701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4373_ clknet_leaf_3_wb_clk_i _0758_ _0356_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3360__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3324_ _1681_ _1698_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__and2_2
XFILLER_0_42_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3255_ _0813_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ net192 _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3186_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\]
+ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2137_ net133 _0933_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2068_ team_10_WB.instance_to_wrap.dispFSM.guesses\[44\] net115 net140 net799 vssd1
+ vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4563__374 vssd1 vssd1 vccd1 vccd1 _4563__374/HI net374 sky130_fd_sc_hd__conb_1
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2191__A team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4709_ net477 vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
XFILLER_0_60_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3351__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2917__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3342__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output66_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3040_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] _1514_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[56\] sky130_fd_sc_hd__mux2_1
XFILLER_0_65_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4547__358 vssd1 vssd1 vccd1 vccd1 _4547__358/HI net358 sky130_fd_sc_hd__conb_1
XFILLER_0_4_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3942_ net242 vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3873_ net260 vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ _1418_ _1426_ _1407_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2755_ net851 _1374_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2686_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\]
+ _1332_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4425_ clknet_leaf_24_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[22\]
+ _0408_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3333__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4356_ clknet_leaf_31_wb_clk_i net756 _0345_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ clknet_leaf_30_wb_clk_i _0677_ _0276_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3238_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ _1638_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3169_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1551_ _1595_ vssd1 vssd1 vccd1
+ vccd1 _0500_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4652__420 vssd1 vssd1 vccd1 vccd1 _4652__420/HI net420 sky130_fd_sc_hd__conb_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4576__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3088__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2540_ _0818_ _0842_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2471_ net613 net128 _1194_ _1209_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4210_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[72\]
+ _0199_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[72\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4141_ clknet_leaf_17_wb_clk_i _0612_ _0140_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4072_ clknet_leaf_36_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[3\]
+ _0092_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3023_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3925_ net270 vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3856_ net287 vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2807_ _1413_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3787_ net272 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2738_ team_10_WB.instance_to_wrap.clock_div.count\[13\] team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ _1362_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout302_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4636__404 vssd1 vssd1 vccd1 vccd1 _4636__404/HI net404 sky130_fd_sc_hd__conb_1
XFILLER_0_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2669_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] _1321_ _1319_ vssd1
+ vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4408_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[5\]
+ _0391_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout212 team_10_WB.instance_to_wrap.gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1
+ net212 sky130_fd_sc_hd__buf_4
Xfanout223 team_10_WB.instance_to_wrap.host_col\[1\] vssd1 vssd1 vccd1 vccd1 net223
+ sky130_fd_sc_hd__buf_2
Xfanout234 net298 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
X_4339_ clknet_leaf_13_wb_clk_i _0729_ _0328_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[62\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_4
Xfanout267 net274 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_4
XFILLER_0_103_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 net281 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_4
XFILLER_0_138_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout289 net296 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2045__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1971_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3710_ net231 vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__inv_2
X_4690_ net458 vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_2
XFILLER_0_43_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3641_ net264 vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3572_ net284 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2744__B1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2523_ net642 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1
+ vccd1 vccd1 _0522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2454_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] net183 vssd1 vssd1 vccd1
+ vccd1 _1200_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2385_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4124_ clknet_leaf_17_wb_clk_i _0595_ _0123_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput1 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
X_4055_ clknet_leaf_7_wb_clk_i _0540_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3006_ team_10_WB.instance_to_wrap.gamelogic.letter\[7\] net125 _1496_ net849 net157
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[39\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4092__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout252_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3908_ net265 vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3839_ net241 vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3295__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4004__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3160__B1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2170_ _0961_ _0960_ _0959_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3099__B net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4742_ net510 vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_2
XFILLER_0_84_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1954_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net147 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4673_ net441 vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_2
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1885_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 _0809_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3624_ net250 vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3555_ net231 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2506_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__or4_1
XANTENNA__3390__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3486_ _1409_ _1436_ _1438_ _1405_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2437_ net608 net131 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2368_ _1091_ _1137_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4748__516 vssd1 vssd1 vccd1 vccd1 _4748__516/HI net516 sky130_fd_sc_hd__conb_1
X_4107_ clknet_leaf_10_wb_clk_i _0578_ _0106_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2299_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4038_ clknet_leaf_35_wb_clk_i _0523_ _0079_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3445__A1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_50 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_61 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_72 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_83 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_94 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input28_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2239__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3436__A1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1998__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold309 team_10_WB.instance_to_wrap.clock_div.count\[19\] vssd1 vssd1 vccd1 vccd1
+ net861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3372__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_3340_ _1694_ _1718_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__nor2_4
XFILLER_0_21_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3271_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ vssd1 vssd1 vccd1 vccd1
+ _1661_ sky130_fd_sc_hd__and4_1
X_2222_ net180 vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__inv_2
XANTENNA__2478__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2153_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2084_ team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] net115 net138 net842 vssd1
+ vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1925__B1_N net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2986_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] net162 _1491_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[24\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2938__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4725_ net493 vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
X_1937_ _0842_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3049__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4656_ net424 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_31_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1868_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1 vccd1 vccd1
+ _0793_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3607_ net261 vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4587_ net63 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3538_ net231 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2189__A team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3469_ team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] net179 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[71\]
+ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2469__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2929__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3354__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2093__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2840_ _1405_ _1426_ _1437_ _1410_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2771_ net858 _1384_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4510_ net321 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4441_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[38\]
+ _0424_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ sky130_fd_sc_hd__dfstp_1
Xhold106 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[21\] vssd1 vssd1
+ vccd1 vccd1 net658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 team_10_WB.instance_to_wrap.host_row1\[72\] vssd1 vssd1 vccd1 vccd1 net669
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold128 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\] vssd1 vssd1 vccd1
+ vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] vssd1 vssd1 vccd1 vccd1
+ net691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4372_ clknet_leaf_23_wb_clk_i _0757_ _0355_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_81_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3323_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ _1698_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__and3_4
XFILLER_0_61_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3254_ net776 _1609_ _1650_ net227 vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__o211a_1
X_2205_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] vssd1 vssd1 vccd1 vccd1 _0993_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3185_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _1608_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710__478 vssd1 vssd1 vccd1 vccd1 _4710__478/HI net478 sky130_fd_sc_hd__conb_1
X_2136_ net213 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0933_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2067_ team_10_WB.instance_to_wrap.dispFSM.guesses\[53\] net141 net107 net673 vssd1
+ vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2191__B team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2969_ net208 net125 _1482_ net782 net157 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[15\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4708_ net476 vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
XFILLER_0_115_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4639_ net407 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3336__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3941_ net250 vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3872_ net251 vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2823_ _0514_ _0513_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2754_ _1373_ _1374_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[19\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4049__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2685_ _1334_ _1335_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[8\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4424_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[21\]
+ _0407_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4355_ clknet_leaf_13_wb_clk_i _0745_ _0344_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[78\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4286_ clknet_leaf_31_wb_clk_i _0676_ _0275_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_96_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3237_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ _1637_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] vssd1 vssd1 vccd1 vccd1
+ _1641_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4530__341 vssd1 vssd1 vccd1 vccd1 _4530__341/HI net341 sky130_fd_sc_hd__conb_1
X_3168_ _1586_ _1590_ _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4569__540 vssd1 vssd1 vccd1 vccd1 net540 _4569__540/LO sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2119_ _0920_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__nor2_2
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3099_ _0789_ net205 vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3254__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3012__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2470_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] net195 team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ net125 vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2523__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4140_ clknet_leaf_18_wb_clk_i _0611_ _0139_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4514__325 vssd1 vssd1 vccd1 vccd1 _4514__325/HI net325 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4071_ clknet_leaf_36_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[2\]
+ _0091_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3022_ net634 net183 _1505_ net200 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[47\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3484__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3924_ net262 vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3855_ net283 vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3846__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2806_ net228 _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3786_ net290 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout128_A _1184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4601__375 vssd1 vssd1 vccd1 vccd1 _4601__375/HI net375 sky130_fd_sc_hd__conb_1
X_2737_ team_10_WB.instance_to_wrap.clock_div.count\[13\] _1362_ net681 vssd1 vssd1
+ vccd1 vccd1 _1363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4675__443 vssd1 vssd1 vccd1 vccd1 _4675__443/HI net443 sky130_fd_sc_hd__conb_1
XFILLER_0_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3057__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2668_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] _1321_ vssd1 vssd1
+ vccd1 vccd1 _1324_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4407_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[4\]
+ _0390_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2599_ _0903_ _1280_ _1282_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__and3b_1
XFILLER_0_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout202 team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 net202
+ sky130_fd_sc_hd__buf_2
Xfanout213 team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1
+ net213 sky130_fd_sc_hd__buf_4
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4716__484 vssd1 vssd1 vccd1 vccd1 _4716__484/HI net484 sky130_fd_sc_hd__conb_1
Xfanout224 _0897_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
Xfanout235 net238 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_4
X_4338_ clknet_leaf_27_wb_clk_i net690 _0327_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout246 net266 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input2_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 net266 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
Xfanout268 net274 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
Xfanout279 net281 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_4
X_4269_ clknet_leaf_50_wb_clk_i _0659_ _0258_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4587__A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_140 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1970_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] net144 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2441__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3640_ net269 vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2992__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4659__427 vssd1 vssd1 vccd1 vccd1 _4659__427/HI net427 sky130_fd_sc_hd__conb_1
XFILLER_0_10_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3571_ net245 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2522_ net579 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1
+ vccd1 vccd1 _0523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2453_ net650 net129 _1185_ _1199_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2384_ _1154_ _1155_ _1087_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4123_ clknet_leaf_24_wb_clk_i _0594_ _0122_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4054_ clknet_leaf_6_wb_clk_i _0539_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput2 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_4
X_3005_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\] net164 _1497_ net832
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[38\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3472__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout245_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3907_ net270 vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3838_ net241 vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3769_ net284 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2196__C1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3160__A1 _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3463__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2974__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3151__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3454__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4780__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4741_ net509 vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_2
XFILLER_0_90_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1953_ net144 net158 vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2965__B2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4672_ net440 vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1884_ team_10_WB.instance_to_wrap.message_reg.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _0808_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3623_ net245 vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3554_ net231 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2505_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[1\] vssd1 vssd1 vccd1 vccd1 _1222_
+ sky130_fd_sc_hd__and3b_1
X_3485_ net588 _1284_ net193 vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2436_ _1193_ _1194_ net639 net129 vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a2bb2o_1
X_2367_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] _1084_ _1140_
+ _1142_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout195_A _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4106_ clknet_leaf_28_wb_clk_i _0577_ _0105_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_2298_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _0823_ _1069_ vssd1 vssd1
+ vccd1 vccd1 _1077_ sky130_fd_sc_hd__nand3_1
XFILLER_0_135_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4037_ clknet_leaf_32_wb_clk_i _0522_ _0078_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3070__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4607__381 vssd1 vssd1 vccd1 vccd1 _4607__381/HI net381 sky130_fd_sc_hd__conb_1
XFILLER_0_1_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_40 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_62 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_73 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_84 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_95 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3381__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3133__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__A2 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1998__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3270_ net294 _1659_ _1660_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__nor3_1
X_2221_ _1001_ _1002_ _1003_ _1006_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__or4_1
XANTENNA__4775__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2883__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2152_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2083_ net685 net141 net107 net716 vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1989__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2985_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__inv_2
XANTENNA__2938__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3060__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4724_ net492 vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1936_ net226 _0857_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__or3b_2
XFILLER_0_44_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4655_ net423 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_114_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1867_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] vssd1 vssd1 vccd1 vccd1
+ _0792_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3606_ net264 vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout110_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4586_ net198 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout208_A team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3537_ net231 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3065__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3468_ net70 net175 _1841_ net227 vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__o211a_1
XANTENNA__2189__B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3115__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2419_ net205 _0942_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__and2_1
X_3399_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] _1688_ _1679_ net206
+ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__o211a_1
XANTENNA__2874__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2636__C _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3051__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input40_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3409__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2770_ _1383_ _1384_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[25\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4440_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[37\]
+ _0423_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold107 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\] vssd1 vssd1 vccd1
+ vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold118 team_10_WB.instance_to_wrap.host_row1\[75\] vssd1 vssd1 vccd1 vccd1 net670
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold129 team_10_WB.instance_to_wrap.clock_div.count\[14\] vssd1 vssd1 vccd1 vccd1
+ net681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4371_ clknet_leaf_23_wb_clk_i _0756_ _0354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3322_ _1683_ _1694_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3253_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] _1607_ _1609_ vssd1 vssd1
+ vccd1 vccd1 _1650_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_47_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2204_ _0946_ net192 _0990_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__o21ai_1
X_3184_ _1603_ _1604_ _1605_ _1606_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ net133 _0932_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2066_ team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] net114 net138 net750 vssd1
+ vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3849__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout158_A _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2472__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3033__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2968_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] net161 _1483_ net209
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[14\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4707_ net475 vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
X_1919_ net222 net223 team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1
+ vccd1 _0842_ sky130_fd_sc_hd__or3_2
XFILLER_0_60_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2899_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\] net152 net123 net714
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[4\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4638_ net406 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ net540 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_64_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3940_ net263 vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3871_ net251 vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
X_4627__395 vssd1 vssd1 vccd1 vccd1 _4627__395/HI net395 sky130_fd_sc_hd__conb_1
XFILLER_0_89_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2822_ net288 _1417_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2753_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[19\]
+ team_10_WB.instance_to_wrap.clock_div.count\[18\] _1367_ vssd1 vssd1 vccd1 vccd1
+ _1374_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2684_ net850 _1332_ _1318_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4423_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[20\]
+ _0406_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_48_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4354_ clknet_leaf_32_wb_clk_i _0744_ _0343_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3305_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__and2b_2
X_4285_ clknet_leaf_13_wb_clk_i _0675_ _0274_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_3236_ net753 _1638_ _1640_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3167_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1278_ _1568_ _1593_ vssd1 vssd1
+ vccd1 vccd1 _1594_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2118_ team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] team_10_WB.instance_to_wrap.buffer.temp_guess\[6\]
+ team_10_WB.instance_to_wrap.buffer.temp_guess\[5\] team_10_WB.instance_to_wrap.buffer.temp_guess\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3098_ net195 net680 net183 _1543_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[85\]
+ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2049_ team_10_WB.instance_to_wrap.dispFSM.guesses\[71\] net142 net108 net722 vssd1
+ vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3088__A3 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3489__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output71_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4553__364 vssd1 vssd1 vccd1 vccd1 _4553__364/HI net364 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4070_ clknet_leaf_36_wb_clk_i net586 _0090_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3021_ _0796_ net183 vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4783__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2039__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4016__CLK clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3923_ net270 vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3854_ net283 vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2805_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[1\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3785_ net289 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2736_ net692 _1362_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[13\]
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2667_ _1318_ _1322_ _1323_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4406_ clknet_leaf_17_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[3\]
+ _0389_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_121_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2598_ _1275_ _1278_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__or2_1
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_4
Xfanout214 team_10_WB.instance_to_wrap.gamelogic.state\[1\] vssd1 vssd1 vccd1 vccd1
+ net214 sky130_fd_sc_hd__buf_2
X_4337_ clknet_leaf_13_wb_clk_i _0727_ _0326_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[60\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _0897_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_1
XANTENNA__3073__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 net238 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_4
Xfanout247 net251 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_4
Xfanout258 net259 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_4
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_4
XFILLER_0_138_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2197__B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4268_ clknet_leaf_0_wb_clk_i _0658_ _0257_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3219_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ net170 vssd1
+ vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3475__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4199_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[61\]
+ _0188_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[61\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4496__307 vssd1 vssd1 vccd1 vccd1 _4496__307/HI net307 sky130_fd_sc_hd__conb_1
XFILLER_0_134_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4537__348 vssd1 vssd1 vccd1 vccd1 _4537__348/HI net348 sky130_fd_sc_hd__conb_1
XFILLER_0_103_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold290 team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] vssd1 vssd1 vccd1 vccd1
+ net842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_130 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_141 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4698__466 vssd1 vssd1 vccd1 vccd1 _4698__466/HI net466 sky130_fd_sc_hd__conb_1
XANTENNA__2729__C1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3570_ net245 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2521_ net565 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] vssd1 vssd1
+ vccd1 vccd1 _0524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1952__B1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2452_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] net183 vssd1 vssd1 vccd1
+ vccd1 _1199_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2383_ _1123_ _1127_ _1136_ _0871_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o31a_1
XFILLER_0_23_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4122_ clknet_leaf_28_wb_clk_i _0593_ _0121_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4053_ clknet_leaf_6_wb_clk_i _0538_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput3 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3004_ _1484_ _1496_ _1497_ _1493_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[37\]
+ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4642__410 vssd1 vssd1 vccd1 vccd1 _4642__410/HI net410 sky130_fd_sc_hd__conb_1
XFILLER_0_8_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3906_ net262 vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout140_A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout238_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3837_ net247 vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2480__B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3068__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3768_ net291 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2719_ _1351_ _1352_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3699_ net240 vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3448__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2974__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3384__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3439__A0 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4740_ net508 vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_2
XFILLER_0_127_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1952_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0874_ net158 _0863_ vssd1
+ vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4671_ net439 vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_2
XFILLER_0_28_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1883_ team_10_WB.instance_to_wrap.message_reg.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _0807_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3622_ net245 vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3553_ net275 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4559__370 vssd1 vssd1 vccd1 vccd1 _4559__370/HI net370 sky130_fd_sc_hd__conb_1
XFILLER_0_84_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2504_ net220 _1221_ _1217_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3484_ net71 net176 _1856_ net227 vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2435_ net130 _1190_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2366_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4105_ clknet_leaf_16_wb_clk_i _0576_ _0104_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2297_ _1069_ _1074_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4036_ clknet_leaf_31_wb_clk_i _0521_ _0077_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2503__A_N net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_52 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_63 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_74 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_85 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_96 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3372__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2220_ net32 net31 _1004_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__or4_1
X_2151_ net164 _0918_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2082_ team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] net114 net138 net864 vssd1
+ vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2984_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] _1191_ _1489_ _1490_
+ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__nand4_4
XFILLER_0_5_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4723_ net491 vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_0_44_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2938__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1935_ _0847_ net194 vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__nand2_2
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4654_ net422 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_47_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1866_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1
+ _0791_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3605_ net249 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4585_ net198 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4754__522 vssd1 vssd1 vccd1 vccd1 _4754__522/HI net522 sky130_fd_sc_hd__conb_1
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3536_ net239 vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3467_ _1704_ _1839_ _1840_ _1838_ _1403_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2418_ _1178_ _1179_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__nor2_1
X_3398_ team_10_WB.instance_to_wrap.host_row2\[43\] team_10_WB.instance_to_wrap.dispFSM.guesses\[19\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2349_ _1122_ _1102_ _1117_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__and3b_1
XANTENNA__3081__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4019_ clknet_leaf_44_wb_clk_i _0504_ _0066_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.unlocked
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4761__526 vssd1 vssd1 vccd1 vccd1 _4761__526/HI net526 sky130_fd_sc_hd__conb_1
XFILLER_0_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2929__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3354__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3780__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input33_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4738__506 vssd1 vssd1 vccd1 vccd1 _4738__506/HI net506 sky130_fd_sc_hd__conb_1
XFILLER_0_41_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold108 team_10_WB.instance_to_wrap.clock_div.count\[27\] vssd1 vssd1 vccd1 vccd1
+ net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] vssd1 vssd1 vccd1
+ vccd1 net671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4370_ clknet_leaf_25_wb_clk_i _0755_ _0353_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3321_ _1686_ _1695_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__and2_2
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3690__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3252_ _1610_ _1649_ net293 vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1922__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2203_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.correct\[0\]
+ team_10_WB.instance_to_wrap.correct\[2\] vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__and3b_2
X_3183_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2134_ net212 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0932_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2065_ team_10_WB.instance_to_wrap.dispFSM.guesses\[55\] net141 net108 net699 vssd1
+ vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__2084__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2967_ _1479_ _1483_ _1484_ _1482_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[13\]
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_91_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4706_ net474 vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
XFILLER_0_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1918_ team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2898_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\] net151 net122 net711
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[3\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_115_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4637_ net405 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_114_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3336__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4568_ net539 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_130_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3519_ net230 vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__inv_2
X_4499_ net310 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4592__551 vssd1 vssd1 vccd1 vccd1 net551 _4592__551/LO sky130_fd_sc_hd__conb_1
XFILLER_0_43_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3870_ net249 vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2821_ _1405_ _1424_ _1425_ _1411_ _1419_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3685__A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2752_ net861 _1372_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2683_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] _1332_ vssd1 vssd1
+ vccd1 vccd1 _1334_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4422_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[19\]
+ _0405_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4353_ clknet_leaf_15_wb_clk_i _0743_ _0342_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[76\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_26_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3304_ _0815_ net206 _1679_ _1681_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4284_ clknet_leaf_30_wb_clk_i net578 _0273_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3235_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\] _1638_ net170 vssd1
+ vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4095__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3166_ _0891_ _0899_ _0906_ net225 vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2117_ team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] team_10_WB.instance_to_wrap.buffer.temp_guess\[2\]
+ team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__or4_1
XFILLER_0_136_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3097_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] net200 vssd1 vssd1 vccd1
+ vccd1 _1543_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2048_ team_10_WB.instance_to_wrap.dispFSM.guesses\[64\] net113 net137 net781 vssd1
+ vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3006__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3999_ clknet_leaf_40_wb_clk_i net553 net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2703__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2004__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4700__468 vssd1 vssd1 vccd1 vccd1 _4700__468/HI net468 sky130_fd_sc_hd__conb_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output64_A net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3020_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\] net184 _1504_ net205
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[46\] sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3484__A1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3922_ net256 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3853_ net242 vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2804_ _1405_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3784_ net291 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2735_ _1361_ _1362_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2666_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1323_ sky130_fd_sc_hd__a21o_1
X_4405_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[2\]
+ _0388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_125_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2597_ _1275_ _1278_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4336_ clknet_leaf_29_wb_clk_i _0726_ _0325_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[59\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout204 net205 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout215 team_10_WB.instance_to_wrap.gamelogic.state\[0\] vssd1 vssd1 vccd1 vccd1
+ net215 sky130_fd_sc_hd__buf_2
Xfanout226 _0846_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout248 net251 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_4
Xfanout259 net265 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_4
X_4267_ clknet_leaf_0_wb_clk_i _0657_ _0256_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3218_ net733 _1626_ _1629_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4198_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[60\]
+ _0187_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[60\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3149_ _0903_ _1277_ _1280_ _1578_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__and4b_1
XFILLER_0_77_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1923__B1_N net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3948__SET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold280 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1
+ net832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold291 team_10_WB.instance_to_wrap.clock_div.count\[23\] vssd1 vssd1 vccd1 vccd1
+ net843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_120 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_131 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_142 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2441__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4520__331 vssd1 vssd1 vccd1 vccd1 _4520__331/HI net331 sky130_fd_sc_hd__conb_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2520_ net570 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1
+ vccd1 vccd1 _0525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1952__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2451_ net640 net132 _1185_ _1198_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2382_ _1123_ _1136_ _1127_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2901__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4121_ clknet_leaf_28_wb_clk_i _0592_ _0120_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4052_ clknet_leaf_6_wb_clk_i _0537_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
X_3003_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\] net159 _1497_ net560
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[36\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_1202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3905_ net258 vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3836_ net262 vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4722__490 vssd1 vssd1 vccd1 vccd1 _4722__490/HI net490 sky130_fd_sc_hd__conb_1
XFILLER_0_7_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3767_ net280 vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3393__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout300_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2718_ net584 _1349_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3698_ net239 vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2649_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__or4bb_1
XANTENNA__3084__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4319_ clknet_leaf_30_wb_clk_i _0709_ _0308_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_138_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4504__315 vssd1 vssd1 vccd1 vccd1 _4504__315/HI net315 sky130_fd_sc_hd__conb_1
XFILLER_0_136_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4771__528 vssd1 vssd1 vccd1 vccd1 _4771__528/HI net528 sky130_fd_sc_hd__conb_1
XFILLER_0_81_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3007__B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4665__433 vssd1 vssd1 vccd1 vccd1 _4665__433/HI net433 sky130_fd_sc_hd__conb_1
XFILLER_0_92_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1951_ team_10_WB.instance_to_wrap.host_message_reg.Cstate team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] _0861_ vssd1 vssd1 vccd1 vccd1
+ _0874_ sky130_fd_sc_hd__nor4_4
X_4706__474 vssd1 vssd1 vccd1 vccd1 _4706__474/HI net474 sky130_fd_sc_hd__conb_1
XFILLER_0_17_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4670_ net438 vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_2
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1882_ team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3621_ net236 vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3375__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3552_ net275 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1925__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2503_ net220 _0889_ net219 vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__and3b_1
XFILLER_0_84_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3483_ _1847_ _1853_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2434_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] _1192_ vssd1 vssd1 vccd1
+ vccd1 _1193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2365_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _0823_ _1069_ _1085_
+ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ clknet_leaf_40_wb_clk_i _0575_ _0103_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2296_ _0841_ _1069_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__or2_2
XFILLER_0_100_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4035_ clknet_leaf_31_wb_clk_i _0520_ _0076_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout250_A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3079__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_20 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_42 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3819_ net250 vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_86 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_97 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3366__B1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2012__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4649__417 vssd1 vssd1 vccd1 vccd1 _4649__417/HI net417 sky130_fd_sc_hd__conb_1
XFILLER_0_138_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3357__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3018__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2150_ net164 _0918_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nor2_1
X_2081_ team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] net142 net108 net703 vssd1
+ vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3688__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2983_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\]
+ _0836_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net160 vssd1 vssd1 vccd1
+ vccd1 _1490_ sky130_fd_sc_hd__a41o_1
XFILLER_0_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4722_ net490 vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
XFILLER_0_5_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1934_ _0843_ net194 vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4653_ net421 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1865_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\] vssd1 vssd1 vccd1 vccd1
+ _0790_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput40 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
X_3604_ net260 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4584_ net197 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3535_ net239 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3466_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1686_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ net207 vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2417_ _1164_ _1167_ _1168_ _1169_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3397_ team_10_WB.instance_to_wrap.host_row1\[59\] _1704_ _1768_ _1773_ vssd1 vssd1
+ vccd1 vccd1 _1774_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2348_ _1102_ _1117_ _1122_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__and3b_1
XFILLER_0_100_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2279_ _0917_ _0948_ _1034_ _1047_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_58_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4018_ clknet_leaf_38_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[2\]
+ net268 vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2007__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4620__391 vssd1 vssd1 vccd1 vccd1 _4620__391/HI net391 sky130_fd_sc_hd__conb_1
XFILLER_0_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold109 team_10_WB.instance_to_wrap.host_row1\[78\] vssd1 vssd1 vccd1 vccd1 net661
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3320_ team_10_WB.instance_to_wrap.host_row2\[40\] net172 _1699_ team_10_WB.instance_to_wrap.host_row1\[48\]
+ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3251_ _1609_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2202_ _0918_ _0972_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3182_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 _1605_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4156__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2133_ _0919_ _0931_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2069__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2064_ team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] net112 net137 net844 vssd1
+ vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2966_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] _1192_ vssd1 vssd1 vccd1
+ vccd1 _1484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4705_ net473 vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
X_1917_ team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__and2b_1
X_2897_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\] net151 net122 net717
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[2\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3149__A_N _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4636_ net404 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_103_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4567_ net538 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3518_ net230 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__inv_2
X_4498_ net309 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3449_ _1821_ _1822_ _1823_ net302 vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__o31a_1
XFILLER_0_99_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2960__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3015__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2820_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2751_ _1371_ _1372_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[18\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2682_ _1318_ _1331_ _1333_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[7\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4421_ clknet_leaf_24_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[18\]
+ _0404_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_125_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2526__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4352_ clknet_leaf_28_wb_clk_i _0742_ _0341_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[75\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3303_ _1680_ _1683_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__nor2_1
X_4283_ clknet_leaf_13_wb_clk_i _0673_ _0272_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_96_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3234_ net665 _1637_ _1639_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3165_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] _1551_ _1591_ _1592_ vssd1 vssd1
+ vccd1 vccd1 _0499_ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2116_ net158 _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__or2_1
X_3096_ net203 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] net189 _1542_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[84\] sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ team_10_WB.instance_to_wrap.dispFSM.guesses\[65\] net109 net135 net848 vssd1
+ vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout163_A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3006__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ clknet_leaf_33_wb_clk_i net555 net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2949_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] net163 _1478_ net213 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[1\] sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1973__C1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4619_ net390 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_108_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2004__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4007__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2453__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3921_ net255 vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2444__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3696__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3852_ net256 vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2803_ _1407_ _0517_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3783_ net280 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2734_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] _1356_ vssd1 vssd1 vccd1 vccd1
+ _1362_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2665_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4404_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[1\]
+ _0387_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_100_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2596_ _1276_ _1280_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__nand2_1
XANTENNA__4062__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4335_ clknet_leaf_29_wb_clk_i _0725_ _0324_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[58\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout205 team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 net205
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout216 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\] vssd1 vssd1 vccd1
+ vccd1 net216 sky130_fd_sc_hd__clkbuf_4
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout238 net243 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
Xfanout249 net251 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_4
X_4266_ clknet_leaf_0_wb_clk_i _0656_ _0255_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3217_ net170 _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3475__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4197_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[59\]
+ _0186_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[59\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3148_ _1571_ _1577_ _1560_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3079_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3350__C_N net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2986__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1961__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\] vssd1 vssd1 vccd1
+ vccd1 net822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\] vssd1 vssd1 vccd1
+ vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold292 team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] vssd1 vssd1 vccd1 vccd1
+ net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_110 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_121 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_132 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2977__B2 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2450_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\] net184 vssd1 vssd1 vccd1
+ vccd1 _1198_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2381_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] _1084_ _1141_
+ _1153_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4120_ clknet_leaf_27_wb_clk_i net600 _0119_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4051_ clknet_leaf_6_wb_clk_i _0536_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3457__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 gpio_in[28] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3002_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\] net159 _1497_ net862
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[35\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3904_ net263 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__inv_2
XANTENNA__2968__B2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3835_ net247 vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3766_ net289 vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2717_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ team_10_WB.instance_to_wrap.clock_div.count\[6\] _1347_ vssd1 vssd1 vccd1 vccd1
+ _1351_ sky130_fd_sc_hd__and4_1
XFILLER_0_131_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3697_ net232 vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__inv_2
XANTENNA__3365__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2648_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[1\] vssd1 vssd1 vccd1 vccd1 _1310_
+ sky130_fd_sc_hd__or3b_2
XFILLER_0_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2579_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] _1259_ _0904_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4318_ clknet_leaf_30_wb_clk_i _0708_ _0307_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[41\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4249_ clknet_leaf_52_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[5\]
+ _0238_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3448__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3081__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4543__354 vssd1 vssd1 vccd1 vccd1 _4543__354/HI net354 sky130_fd_sc_hd__conb_1
XFILLER_0_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3384__A1 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3136__A1 _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2895__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1950_ _0841_ _0871_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__or2_2
XFILLER_0_84_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1881_ team_10_WB.instance_to_wrap.gamelogic.green vssd1 vssd1 vccd1 vccd1 _0806_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3620_ net244 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3551_ net279 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1925__A2 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2502_ net219 _1220_ _1217_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3482_ _1727_ _1854_ _1403_ _1689_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2433_ net661 net131 _1191_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2364_ _1138_ _1139_ _1088_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__o21a_1
X_4103_ clknet_leaf_40_wb_clk_i _0574_ _0102_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2295_ _0840_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4034_ clknet_leaf_31_wb_clk_i _0519_ _0075_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4527__338 vssd1 vssd1 vccd1 vccd1 _4527__338/HI net338 sky130_fd_sc_hd__conb_1
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout243_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_21 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_54 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3818_ net259 vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__inv_2
XANTENNA_65 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_76 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_87 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_98 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3749_ net278 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2012__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2877__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4688__456 vssd1 vssd1 vccd1 vccd1 _4688__456/HI net456 sky130_fd_sc_hd__conb_1
XFILLER_0_138_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2644__A3 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4729__497 vssd1 vssd1 vccd1 vccd1 _4729__497/HI net497 sky130_fd_sc_hd__conb_1
XFILLER_0_69_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3357__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4632__400 vssd1 vssd1 vccd1 vccd1 _4632__400/HI net400 sky130_fd_sc_hd__conb_1
XFILLER_0_123_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2080_ team_10_WB.instance_to_wrap.dispFSM.guesses\[32\] net113 net137 net758 vssd1
+ vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2979__A1_N _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2982_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] _0837_ net160 vssd1 vssd1 vccd1
+ vccd1 _1489_ sky130_fd_sc_hd__a41o_1
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4721_ net489 vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
X_1933_ _0850_ net194 vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4652_ net420 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1864_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1 vccd1 vccd1
+ _0789_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput30 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3603_ net269 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput41 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
X_4583_ net546 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_0_12_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3534_ net237 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3465_ team_10_WB.instance_to_wrap.host_row1\[62\] team_10_WB.instance_to_wrap.dispFSM.msg\[6\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__mux2_1
X_2416_ _1177_ net229 _0849_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__and3b_2
X_3396_ team_10_WB.instance_to_wrap.host_row1\[43\] _1693_ _1770_ _1771_ _1772_ vssd1
+ vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__a2111o_1
X_2347_ _1117_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2278_ _0950_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4017_ clknet_leaf_34_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[1\]
+ net276 vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3036__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input19_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4549__360 vssd1 vssd1 vccd1 vccd1 _4549__360/HI net360 sky130_fd_sc_hd__conb_1
XFILLER_0_98_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3250_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\] _1608_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2201_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] _0989_ _0973_ vssd1
+ vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o21a_1
X_3181_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__or4b_1
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2132_ net211 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2063_ team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] net109 net134 net775 vssd1
+ vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2965_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\] net161 _1483_ net210
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[12\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__1947__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4704_ net472 vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XFILLER_0_127_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1916_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\] vssd1 vssd1 vccd1 vccd1
+ _0839_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2896_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\] net153 _1473_ net713
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[1\]
+ sky130_fd_sc_hd__o22a_1
X_4635_ net403 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ net537 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_114_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3517_ net230 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__inv_2
X_4497_ net308 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3448_ team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] net169 net167 team_10_WB.instance_to_wrap.dispFSM.msg\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3379_ team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] net171 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[2\]
+ _1756_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4744__512 vssd1 vssd1 vccd1 vccd1 _4744__512/HI net512 sky130_fd_sc_hd__conb_1
XFILLER_0_54_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ team_10_WB.instance_to_wrap.clock_div.count\[18\] _1365_ vssd1 vssd1 vccd1 vccd1
+ _1372_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2681_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4420_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[17\]
+ _0403_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_48_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4351_ clknet_leaf_29_wb_clk_i _0741_ _0340_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[74\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _1681_ _1682_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4282_ clknet_leaf_29_wb_clk_i _0672_ _0271_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3233_ net170 _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__nor2_1
X_3164_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] _1278_ _1568_ _0903_ vssd1 vssd1
+ vccd1 vccd1 _1592_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2115_ _0916_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__or2_2
XFILLER_0_136_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3095_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] net196 vssd1 vssd1 vccd1
+ vccd1 _1542_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ team_10_WB.instance_to_wrap.dispFSM.guesses\[66\] net110 net134 net786 vssd1
+ vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout156_A _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3997_ clknet_leaf_42_wb_clk_i _0487_ _0065_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2948_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] net162 _1478_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[0\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2879_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\] vssd1 vssd1 vccd1 vccd1
+ _1463_ sky130_fd_sc_hd__and3b_1
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4203__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[65\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4618_ net389 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_130_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4549_ net360 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_44_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3478__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3469__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3920_ net257 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3851_ net242 vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2802_ _1409_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3782_ net289 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2733_ net814 _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2664_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1321_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4403_ clknet_leaf_16_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[0\]
+ _0386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_125_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2595_ _0908_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4334_ clknet_leaf_30_wb_clk_i _0724_ _0323_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[57\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout206 net207 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
Xfanout228 _0018_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout239 net243 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_4
X_4265_ clknet_leaf_56_wb_clk_i _0655_ _0254_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3216_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] _1626_ vssd1 vssd1 vccd1
+ vccd1 _1628_ sky130_fd_sc_hd__and2_1
X_4196_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[58\]
+ _0185_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[58\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2132__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3147_ _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout273_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3078_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] _1533_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[75\] sky130_fd_sc_hd__mux2_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2029_ net193 _0909_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold260 team_10_WB.instance_to_wrap.dispFSM.guesses\[70\] vssd1 vssd1 vccd1 vccd1
+ net812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] vssd1 vssd1 vccd1 vccd1
+ net823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_10_WB.instance_to_wrap.dispFSM.guesses\[14\] vssd1 vssd1 vccd1 vccd1
+ net834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold293 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] vssd1 vssd1 vccd1
+ vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2966__A team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_100 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_111 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_122 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_133 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2206__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2380_ _0871_ _1088_ _1152_ _1075_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2901__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4050_ clknet_leaf_6_wb_clk_i _0535_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3001_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\] net159 _1497_ net558
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[34\]
+ sky130_fd_sc_hd__o22a_1
Xinput6 gpio_in[37] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3903_ net248 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3090__A1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2116__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3834_ net258 vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3765_ net278 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1955__A team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2716_ _1171_ _1349_ _1350_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[5\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__3393__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3696_ net232 vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout119_A _0875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2647_ _1307_ _1308_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2578_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] _0898_ _0901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4317_ clknet_leaf_14_wb_clk_i _0707_ _0306_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[40\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3381__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4248_ clknet_leaf_52_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[4\]
+ _0237_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4179_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[41\]
+ _0168_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[41\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3384__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1880_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1 vccd1
+ _0805_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3550_ net277 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__inv_2
XANTENNA__3375__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2501_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3481_ team_10_WB.instance_to_wrap.host_row2\[71\] team_10_WB.instance_to_wrap.dispFSM.guesses\[47\]
+ net6 vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2432_ net192 _1186_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2363_ net226 _0847_ _0853_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__and3b_1
XANTENNA__2886__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4102_ clknet_leaf_40_wb_clk_i _0573_ _0101_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2294_ _0859_ _0865_ _1071_ _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4033_ clknet_leaf_10_wb_clk_i _0518_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_33 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_44 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_55 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3817_ net259 vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
XANTENNA_66 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_77 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_88 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_99 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3748_ net292 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3679_ net265 vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4510__321 vssd1 vssd1 vccd1 vccd1 _4510__321/HI net321 sky130_fd_sc_hd__conb_1
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3357__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4712__480 vssd1 vssd1 vccd1 vccd1 _4712__480/HI net480 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2981_ net208 _1485_ _1488_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[23\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4720_ net488 vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
X_1932_ team_10_WB.instance_to_wrap.host_col\[3\] net222 team_10_WB.instance_to_wrap.host_col\[1\]
+ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__or4_2
XFILLER_0_51_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4651_ net419 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_127_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1863_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1
+ _0788_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
X_3602_ net288 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__inv_2
Xinput31 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_4582_ net545 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3533_ net246 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3464_ _1828_ _1831_ _1837_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2415_ net229 _1171_ net554 vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3395_ team_10_WB.instance_to_wrap.host_row1\[51\] _1699_ net177 team_10_WB.instance_to_wrap.host_row2\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2346_ _0829_ _1121_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _1122_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2277_ _1054_ _1055_ _1058_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__and3b_1
XFILLER_0_97_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4016_ clknet_3_3_0_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[0\]
+ net268 vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4206__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4655__423 vssd1 vssd1 vccd1 vccd1 _4655__423/HI net423 sky130_fd_sc_hd__conb_1
XFILLER_0_132_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2200_ _0919_ _0971_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3180_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__or4b_1
XFILLER_0_98_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2131_ net133 _0930_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2062_ team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] net110 net134 net783 vssd1
+ vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2069__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2964_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] net160 _1483_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[11\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4703_ net471 vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
X_1915_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] vssd1 vssd1 vccd1 vccd1
+ _0838_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2895_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\] net153 net120 net725
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[0\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4634_ net402 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
X_4639__407 vssd1 vssd1 vccd1 vccd1 _4639__407/HI net407 sky130_fd_sc_hd__conb_1
XFILLER_0_128_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4565_ net536 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3516_ net230 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__inv_2
X_4496_ net307 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_106_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3447_ team_10_WB.instance_to_wrap.dispFSM.guesses\[21\] net172 net166 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\]
+ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3378_ team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] _1715_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[66\]
+ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2329_ _0819_ _0849_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] vssd1
+ vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2018__B net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1873__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input31_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2456__C1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2471__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2680_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ _1327_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4350_ clknet_leaf_31_wb_clk_i _0740_ _0339_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[73\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3301_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net206 vssd1 vssd1 vccd1
+ vccd1 _1682_ sky130_fd_sc_hd__nor2_1
XANTENNA__2931__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4281_ clknet_leaf_13_wb_clk_i _0671_ _0270_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3232_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] _1637_ vssd1 vssd1 vccd1
+ vccd1 _1638_ sky130_fd_sc_hd__and2_1
X_3163_ _1586_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2114_ net215 net214 vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand2_1
X_3094_ net204 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] net188 _1541_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[83\] sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ team_10_WB.instance_to_wrap.dispFSM.guesses\[67\] net111 net136 net816 vssd1
+ vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3996_ clknet_leaf_42_wb_clk_i _0486_ _0064_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout149_A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2947_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] net162 _1475_ _1476_ _1477_
+ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2878_ net191 _1462_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[2\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__1973__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4617_ net388 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4548_ net359 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_130_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2922__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4479_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[36\]
+ _0462_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2029__A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2438__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1868__A team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1964__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1964__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2913__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3850_ net255 vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2801_ net227 _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3781_ net277 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2732_ _1359_ _1360_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[11\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2663_ net651 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\] _1320_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4402_ clknet_leaf_47_wb_clk_i _0787_ _0385_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2594_ _0890_ net225 net220 vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2904__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4333_ clknet_leaf_14_wb_clk_i _0723_ _0322_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[56\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout207 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\] vssd1 vssd1 vccd1
+ vccd1 net207 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout218 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] vssd1 vssd1 vccd1
+ vccd1 net218 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2380__B2 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 _0821_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4264_ clknet_leaf_56_wb_clk_i _0654_ _0253_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3215_ net877 _1624_ _1627_ _1611_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4195_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[57\]
+ _0184_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[57\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3146_ _1573_ _1574_ _1569_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3077_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout266_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2028_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3979_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[16\]
+ _0047_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\] vssd1 vssd1 vccd1 vccd1
+ net802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold261 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\] vssd1 vssd1 vccd1
+ vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold272 team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] vssd1 vssd1 vccd1 vccd1
+ net824 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2371__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold283 team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] vssd1 vssd1 vccd1 vccd1
+ net835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\] vssd1 vssd1 vccd1 vccd1
+ net846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3320__B1 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_101 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_112 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_123 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_134 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2206__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3387__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3000_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\] net159 _1497_ net605
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[33\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput7 wb_rst_i vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4566__537 vssd1 vssd1 vccd1 vccd1 net537 _4566__537/LO sky130_fd_sc_hd__conb_1
XFILLER_0_73_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3902_ net248 vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3833_ net258 vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3378__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3764_ net292 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2715_ team_10_WB.instance_to_wrap.clock_div.count\[4\] _1347_ team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3695_ net232 vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2646_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] _0827_ team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2577_ _1254_ _1255_ _1260_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4316_ clknet_leaf_31_wb_clk_i _0706_ _0305_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4247_ clknet_leaf_51_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[3\]
+ _0236_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4178_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[40\]
+ _0167_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[40\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3129_ _1557_ _1559_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3369__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2895__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4589__548 vssd1 vssd1 vccd1 vccd1 net548 _4589__548/LO sky130_fd_sc_hd__conb_1
XFILLER_0_38_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2500_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\] team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\]
+ net220 net217 vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__or4b_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3480_ team_10_WB.instance_to_wrap.host_row2\[55\] net168 _1848_ _1852_ vssd1 vssd1
+ vccd1 vccd1 _1853_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2431_ net192 _1186_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2362_ _1091_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4101_ clknet_leaf_40_wb_clk_i _0572_ _0100_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2293_ _0843_ net226 net194 _0858_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_58_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4032_ clknet_leaf_9_wb_clk_i _0517_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2127__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3816_ net249 vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout131_A _1183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_56 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_89 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3747_ net272 vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3678_ net258 vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2629_ _0807_ _0808_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.blue sky130_fd_sc_hd__nor2_4
XFILLER_0_41_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1876__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2014__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2980_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] net159 _1488_ team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[22\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1931_ net226 _0848_ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1
+ vccd1 _0854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4650_ net418 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_115_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput10 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_4
X_3601_ net285 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput21 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
X_4581_ net197 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
Xinput32 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput43 wbs_we_i vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3532_ net246 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3463_ team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] net177 _1832_ _1836_ vssd1
+ vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__a211o_1
XANTENNA__2308__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2414_ team_10_WB.instance_to_wrap.clock_div.count\[6\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ _1170_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__or4_4
XFILLER_0_0_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3394_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net206 _1681_ _1686_
+ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2345_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _0870_ _1118_ _1120_
+ _0828_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__a32o_1
X_4533__344 vssd1 vssd1 vccd1 vccd1 _4533__344/HI net344 sky130_fd_sc_hd__conb_1
XFILLER_0_97_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2276_ _0791_ net208 _1050_ _1053_ _1057_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4015_ clknet_leaf_32_wb_clk_i _0503_ net273 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4779_ net531 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_105_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4694__462 vssd1 vssd1 vccd1 vccd1 _4694__462/HI net462 sky130_fd_sc_hd__conb_1
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4042__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2483__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4517__328 vssd1 vssd1 vccd1 vccd1 _4517__328/HI net328 sky130_fd_sc_hd__conb_1
XFILLER_0_24_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2130_ net210 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2061_ team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] net111 net136 net809 vssd1
+ vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3423__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2963_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] net160 _1483_ net212
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[10\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4702_ net470 vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
XFILLER_0_127_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1914_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\] vssd1 vssd1 vccd1 vccd1
+ _0837_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2894_ net158 net149 vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__nand2_2
XFILLER_0_72_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4604__378 vssd1 vssd1 vccd1 vccd1 _4604__378/HI net378 sky130_fd_sc_hd__conb_1
XFILLER_0_127_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4633_ net401 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
X_4678__446 vssd1 vssd1 vccd1 vccd1 _4678__446/HI net446 sky130_fd_sc_hd__conb_1
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4564_ net535 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3515_ net230 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__inv_2
X_4495_ net306 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
X_4719__487 vssd1 vssd1 vccd1 vccd1 _4719__487/HI net487 sky130_fd_sc_hd__conb_1
XFILLER_0_106_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3446_ team_10_WB.instance_to_wrap.dispFSM.guesses\[77\] _1715_ _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[13\]
+ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3377_ team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] net179 net177 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\]
+ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout296_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2701__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2328_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\] _0858_ vssd1 vssd1
+ vccd1 vccd1 _1104_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2259_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0798_ _1036_ _1037_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_34_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1976__C1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1991__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2940__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4088__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3300_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _0817_ vssd1 vssd1 vccd1
+ vccd1 _1681_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4280_ clknet_leaf_14_wb_clk_i _0670_ _0269_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3231_ _1637_ _1611_ _1636_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and3b_1
XFILLER_0_123_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3162_ _0812_ net4 _0906_ _1582_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2113_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__nand2b_1
X_3093_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net196 vssd1 vssd1 vccd1
+ vccd1 _1541_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2044_ team_10_WB.instance_to_wrap.dispFSM.guesses\[68\] net112 net137 net691 vssd1
+ vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3995_ clknet_leaf_42_wb_clk_i _0485_ _0063_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2135__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2946_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\]
+ net160 vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__a41o_1
XANTENNA__3411__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2877_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] _1461_ vssd1 vssd1 vccd1
+ vccd1 _1462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4616_ net387 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XANTENNA_fanout211_A team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4547_ net358 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4539__350 vssd1 vssd1 vccd1 vccd1 _4539__350/HI net350 sky130_fd_sc_hd__conb_1
XFILLER_0_130_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4478_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[35\]
+ _0461_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3429_ net302 team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _0815_ net207 vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__o2111a_1
XANTENNA__3950__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3478__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2438__B1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2989__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4774__529 vssd1 vssd1 vccd1 vccd1 _4774__529/HI net529 sky130_fd_sc_hd__conb_1
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3469__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2429__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2800_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[4\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3780_ net294 vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2731_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ _1356_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2662_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ _1318_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4401_ clknet_leaf_4_wb_clk_i _0786_ _0384_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2593_ _0910_ _1276_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__nand2_2
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_4332_ clknet_leaf_31_wb_clk_i _0722_ _0321_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout208 team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1
+ net208 sky130_fd_sc_hd__buf_4
Xfanout219 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1 vccd1
+ vccd1 net219 sky130_fd_sc_hd__buf_2
X_4263_ clknet_leaf_56_wb_clk_i _0653_ _0252_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3214_ _1626_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4194_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[56\]
+ _0183_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[56\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3145_ _1569_ _1573_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3076_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] _1532_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[74\] sky130_fd_sc_hd__mux2_1
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2027_ _0888_ _0908_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout259_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ clknet_leaf_43_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[15\]
+ _0046_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2929_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] net150 net121 net773
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[34\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4734__502 vssd1 vssd1 vccd1 vccd1 _4734__502/HI net502 sky130_fd_sc_hd__conb_1
XFILLER_0_130_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold240 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] vssd1 vssd1 vccd1
+ vccd1 net792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] vssd1 vssd1 vccd1 vccd1
+ net803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold262 team_10_WB.instance_to_wrap.clock_div.count\[12\] vssd1 vssd1 vccd1 vccd1
+ net814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] vssd1 vssd1 vccd1 vccd1
+ net825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold284 team_10_WB.instance_to_wrap.clock_div.count\[2\] vssd1 vssd1 vccd1 vccd1
+ net836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] vssd1 vssd1 vccd1 vccd1
+ net847 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4617__388 vssd1 vssd1 vccd1 vccd1 _4617__388/HI net388 sky130_fd_sc_hd__conb_1
XFILLER_0_92_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_102 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1879__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_113 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_124 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3084__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_135 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2898__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_4
XFILLER_0_127_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3901_ net250 vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3090__A3 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3832_ net263 vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3763_ net271 vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2714_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ _1347_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3694_ net240 vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2645_ net1 net158 team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1
+ vccd1 vccd1 _1307_ sky130_fd_sc_hd__and3b_1
XFILLER_0_112_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2576_ net217 net224 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] vssd1
+ vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4315_ clknet_leaf_12_wb_clk_i _0705_ _0304_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[38\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_26_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4246_ clknet_leaf_52_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[2\]
+ _0235_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4177_ clknet_leaf_47_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[2\]
+ _0166_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__dfrtp_1
X_3128_ _1286_ _1288_ _1291_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3066__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3059_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4149__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3154__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2032__A1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2430_ _0993_ _1185_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__and2_2
XFILLER_0_62_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2361_ _1096_ _1131_ _1135_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4100_ clknet_leaf_8_wb_clk_i _0571_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2292_ _0842_ _0866_ _1070_ _0865_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4031_ clknet_leaf_9_wb_clk_i _0516_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3296__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2271__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_13 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3815_ net248 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
XANTENNA_35 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_46 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_57 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_68 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3746_ net290 vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3677_ net256 vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2628_ _0009_ _0010_ _0008_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2797__B net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2559_ net215 _0952_ _1024_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4229_ clknet_leaf_56_wb_clk_i _0645_ _0218_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2014__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2500__B team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1930_ net223 _0851_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3600_ net260 vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__inv_2
Xinput11 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_4580_ net198 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput22 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput33 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3531_ net246 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3462_ team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] net169 _1833_ _1835_ vssd1
+ vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2413_ _1167_ _1173_ _1174_ _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3393_ team_10_WB.instance_to_wrap.host_row2\[83\] net171 net165 team_10_WB.instance_to_wrap.host_row2\[75\]
+ _1769_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2344_ _0823_ _1857_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] vssd1 vssd1
+ vccd1 vccd1 _1120_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2275_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] _1056_ vssd1 vssd1
+ vccd1 vccd1 _1057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4014_ clknet_leaf_33_wb_clk_i _0502_ net273 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[6\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2244__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2244__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4778_ net181 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3729_ net252 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold286_A team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2235__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2235__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1994__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_4556__367 vssd1 vssd1 vccd1 vccd1 _4556__367/HI net367 sky130_fd_sc_hd__conb_1
XFILLER_0_123_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2060_ team_10_WB.instance_to_wrap.dispFSM.guesses\[52\] net115 net140 net760 vssd1
+ vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2962_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\] net162 _1483_ net213 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[9\] sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4701_ net469 vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
X_1913_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\] vssd1 vssd1 vccd1 vccd1
+ _0836_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2893_ net163 net155 vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4632_ net400 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_72_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4500__311 vssd1 vssd1 vccd1 vccd1 _4500__311/HI net311 sky130_fd_sc_hd__conb_1
X_4563_ net374 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XFILLER_0_128_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3514_ net235 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2421__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4494_ net305 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_106_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3445_ _0821_ _1819_ _1817_ _1812_ _1807_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3376_ team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] net172 net169 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\]
+ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2327_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\] _0854_ vssd1 vssd1
+ vccd1 vccd1 _1103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout289_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2258_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0798_ _0799_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2189_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] net209 vssd1 vssd1 vccd1
+ vccd1 _0978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3414__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4702__470 vssd1 vssd1 vccd1 vccd1 _4702__470/HI net470 sky130_fd_sc_hd__conb_1
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2940__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2456__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3405__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1967__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2241__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2392__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751__519 vssd1 vssd1 vccd1 vccd1 _4751__519/HI net519 sky130_fd_sc_hd__conb_1
XANTENNA__2931__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3230_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ _1633_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3161_ team_10_WB.instance_to_wrap.dispFSM.msg\[2\] _0886_ _1274_ _1581_ _1589_ vssd1
+ vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__o32a_1
XFILLER_0_59_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2112_ team_10_WB.instance_to_wrap.dispFSM.guesses\[0\] net113 net139 team_10_WB.instance_to_wrap.dispFSM.guesses\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__o22a_1
X_3092_ net203 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] net188 _1540_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[82\] sky130_fd_sc_hd__a31o_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2043_ team_10_WB.instance_to_wrap.dispFSM.guesses\[77\] net141 net107 net727 vssd1
+ vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4645__413 vssd1 vssd1 vccd1 vccd1 _4645__413/HI net413 sky130_fd_sc_hd__conb_1
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3994_ clknet_leaf_42_wb_clk_i _0484_ _0062_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4032__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2945_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] net125 _1474_ vssd1
+ vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1958__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2876_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] net221 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4615_ team_10_WB.instance_to_wrap.gamelogic.red vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2151__A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4546_ net357 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_111_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout204_A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2922__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4477_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[34\]
+ _0460_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3428_ team_10_WB.instance_to_wrap.host_row1\[53\] net301 _1699_ vssd1 vssd1 vccd1
+ vccd1 _1803_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3332__C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3359_ team_10_WB.instance_to_wrap.host_row1\[41\] _1693_ _1703_ team_10_WB.instance_to_wrap.host_row1\[65\]
+ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3710__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600__552 vssd1 vssd1 vccd1 vccd1 net552 _4600__552/LO sky130_fd_sc_hd__conb_1
XFILLER_0_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2913__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2126__A0 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4055__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2730_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ net873 vssd1 vssd1
+ vccd1 vccd1 _1359_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2661_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\] _1319_ vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[0\] sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4400_ clknet_leaf_47_wb_clk_i _0785_ _0383_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\]
+ sky130_fd_sc_hd__dfrtp_4
X_2592_ _0910_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4331_ clknet_leaf_13_wb_clk_i _0721_ _0320_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[54\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout209 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1
+ net209 sky130_fd_sc_hd__clkbuf_4
X_4262_ clknet_leaf_57_wb_clk_i _0652_ _0251_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3213_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\] _1621_ vssd1 vssd1 vccd1 vccd1
+ _1626_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4193_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[55\]
+ _0182_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[55\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3144_ _1557_ _1571_ _1572_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3075_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__mux2_1
XANTENNA__3530__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2026_ _0888_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3977_ clknet_3_0_0_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[14\]
+ _0045_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1985__A team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3396__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2928_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] net149 net120 net780
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[33\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2859_ _1450_ _1451_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold230 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\] vssd1 vssd1 vccd1 vccd1
+ net782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold241 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\] vssd1 vssd1 vccd1
+ vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ net340 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
Xhold252 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] vssd1 vssd1 vccd1
+ vccd1 net804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\] vssd1 vssd1 vccd1
+ vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold274 team_10_WB.instance_to_wrap.clock_div.count\[25\] vssd1 vssd1 vccd1 vccd1
+ net826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] vssd1 vssd1 vccd1 vccd1
+ net837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 team_10_WB.instance_to_wrap.dispFSM.guesses\[73\] vssd1 vssd1 vccd1 vccd1
+ net848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3320__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_103 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_114 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_125 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_136 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3387__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_4
XFILLER_0_86_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ net264 vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3831_ net248 vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3378__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3762_ net294 vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4757__525 vssd1 vssd1 vccd1 vccd1 _4757__525/HI net525 sky130_fd_sc_hd__conb_1
X_2713_ net675 _1347_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
X_3693_ net240 vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2644_ _0923_ _0947_ _1302_ _0924_ _0922_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[3\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_112_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2575_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] net224 net217 vssd1
+ vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__nand3b_1
XANTENNA__2889__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4314_ clknet_leaf_32_wb_clk_i _0704_ _0303_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4245_ clknet_leaf_52_wb_clk_i net652 _0234_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4176_ clknet_leaf_45_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[1\]
+ _0165_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3127_ _1862_ _1555_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] vssd1
+ vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout271_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3058_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _1523_ net199 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[65\] sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2009_ net216 net217 net219 net220 vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__nor4_1
XFILLER_0_93_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3369__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2032__A2 _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2360_ _1124_ _1134_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__xor2_1
X_4572__543 vssd1 vssd1 vccd1 vccd1 net543 _4572__543/LO sky130_fd_sc_hd__conb_1
XFILLER_0_23_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2291_ net5 _0844_ net194 vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4030_ clknet_leaf_9_wb_clk_i _0515_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2099__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_14 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_25 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ net248 vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2424__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_47 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2559__B1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_69 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3745_ net289 vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3676_ net241 vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout117_A _0875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2627_ net875 _1074_ _1297_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2558_ _1243_ _1247_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2489_ net593 net128 _1189_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] vssd1
+ vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__o22a_1
X_4228_ clknet_leaf_56_wb_clk_i _0644_ _0217_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4159_ clknet_leaf_42_wb_clk_i _0628_ _0148_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2014__A2 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2500__C net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2486__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput23 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3530_ net246 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3461_ team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] net179 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[70\]
+ _1834_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2412_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3392_ team_10_WB.instance_to_wrap.host_row1\[75\] _1708_ net178 team_10_WB.instance_to_wrap.host_row2\[59\]
+ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2343_ _0870_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2274_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0800_ _1051_ _1052_ _1049_
+ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__a221o_1
X_4013_ clknet_leaf_33_wb_clk_i _0501_ net268 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2419__A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3441__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2244__A2 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3441__B2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4777_ net530 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3944__RESET_B _0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1989_ net856 net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] vssd1
+ vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3728_ net240 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2952__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3659_ net289 vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3713__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2483__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2235__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1994__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1994__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2459__C1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2474__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3423__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2961_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\] net162 _1483_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[8\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ net468 vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
XFILLER_0_57_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1912_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\] vssd1 vssd1 vccd1 vccd1
+ _0835_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2892_ net191 _1471_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_71_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4631_ net399 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4562_ net373 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_25_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3513_ net235 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2421__B net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4493_ net304 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_106_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3444_ team_10_WB.instance_to_wrap.host_row2\[45\] net172 net167 team_10_WB.instance_to_wrap.host_row1\[61\]
+ _1818_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3375_ team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] net166 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3533__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2162__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2326_ _1100_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2257_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] net213 vssd1 vssd1 vccd1
+ vccd1 _1039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout184_A _0995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2188_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net212 vssd1 vssd1 vccd1
+ vccd1 _0977_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3414__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1976__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3708__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2925__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3162__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2456__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2208__A2 _0995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4523__334 vssd1 vssd1 vccd1 vccd1 _4523__334/HI net334 sky130_fd_sc_hd__conb_1
XFILLER_0_13_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3341__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3160_ _0903_ _1588_ net193 vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2111_ team_10_WB.instance_to_wrap.dispFSM.guesses\[1\] net109 net135 net871 vssd1
+ vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe vssd1 vssd1 vccd1 vccd1
+ net553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3091_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] net196 vssd1 vssd1 vccd1
+ vccd1 _1540_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2042_ team_10_WB.instance_to_wrap.dispFSM.guesses\[70\] net113 net137 net805 vssd1
+ vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4610__384 vssd1 vssd1 vccd1 vccd1 _4610__384/HI net384 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4684__452 vssd1 vssd1 vccd1 vccd1 _4684__452/HI net452 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2416__B net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3993_ clknet_leaf_40_wb_clk_i _0483_ _0061_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4725__493 vssd1 vssd1 vccd1 vccd1 _4725__493/HI net493 sky130_fd_sc_hd__conb_1
XFILLER_0_17_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2944_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] _0831_ net162 vssd1 vssd1
+ vccd1 vccd1 _1475_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2875_ net191 _1460_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[1\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2432__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4614_ team_10_WB.instance_to_wrap.gamelogic.green vssd1 vssd1 vccd1 vccd1 net73
+ sky130_fd_sc_hd__buf_1
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2907__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4545_ net356 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4476_ clknet_leaf_48_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[33\]
+ _0459_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_64_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3427_ team_10_WB.instance_to_wrap.host_row2\[61\] team_10_WB.instance_to_wrap.dispFSM.guesses\[37\]
+ net300 vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3358_ team_10_WB.instance_to_wrap.host_row2\[41\] net172 net171 team_10_WB.instance_to_wrap.host_row2\[81\]
+ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2309_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] _1076_ _1077_
+ net163 vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__a31o_1
X_3289_ _1672_ _1673_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2438__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4507__318 vssd1 vssd1 vccd1 vccd1 _4507__318/HI net318 sky130_fd_sc_hd__conb_1
XFILLER_0_119_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3020__C1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4668__436 vssd1 vssd1 vccd1 vccd1 _4668__436/HI net436 sky130_fd_sc_hd__conb_1
XFILLER_0_95_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2429__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4709__477 vssd1 vssd1 vccd1 vccd1 _4709__477/HI net477 sky130_fd_sc_hd__conb_1
XFILLER_0_86_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2660_ _1307_ _1310_ _1313_ _1317_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_67_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2591_ _0908_ _1219_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ clknet_leaf_27_wb_clk_i _0720_ _0319_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4261_ clknet_leaf_1_wb_clk_i _0651_ _0250_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.red
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3212_ net789 _1622_ _1625_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4192_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[54\]
+ _0181_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[54\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3143_ _1557_ _1572_ _1571_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3811__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3074_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] _1531_ net199 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[73\] sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2025_ net3 _0901_ _0907_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2427__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4582__545 vssd1 vssd1 vccd1 vccd1 net545 _4582__545/LO sky130_fd_sc_hd__conb_1
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3976_ clknet_leaf_43_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[13\]
+ _0044_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2053__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2927_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] net149 net120 net793
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[32\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2858_ net868 _1448_ net174 vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2789_ _1393_ _1395_ _1396_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] vssd1 vssd1 vccd1
+ vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4528_ net339 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_41_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold231 team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] vssd1 vssd1 vccd1 vccd1
+ net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold242 team_10_WB.instance_to_wrap.dispFSM.guesses\[24\] vssd1 vssd1 vccd1 vccd1
+ net794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 team_10_WB.instance_to_wrap.dispFSM.guesses\[78\] vssd1 vssd1 vccd1 vccd1
+ net805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 team_10_WB.instance_to_wrap.dispFSM.guesses\[75\] vssd1 vssd1 vccd1 vccd1
+ net816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 team_10_WB.instance_to_wrap.clock_div.count\[8\] vssd1 vssd1 vccd1 vccd1
+ net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold286 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 net838
+ sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[16\]
+ _0442_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\]
+ sky130_fd_sc_hd__dfstp_1
Xhold297 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\] vssd1 vssd1 vccd1 vccd1
+ net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3721__A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_104 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_115 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_126 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_137 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2898__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4529__340 vssd1 vssd1 vccd1 vccd1 _4529__340/HI net340 sky130_fd_sc_hd__conb_1
XFILLER_0_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3830_ net259 vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3761_ net284 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2712_ _1347_ _1348_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3692_ net279 vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2643_ _0953_ _1306_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2574_ net219 net224 vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4313_ clknet_leaf_12_wb_clk_i _0703_ _0302_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3017__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4244_ clknet_leaf_51_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[0\]
+ _0233_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4175_ clknet_leaf_45_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[0\]
+ _0164_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3126_ _1286_ _1554_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__nor3_2
XFILLER_0_39_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3057_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\]
+ net185 vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout264_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2008_ net219 _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3959_ clknet_leaf_45_wb_clk_i _0010_ _0027_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3716__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4045__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4630__398 vssd1 vssd1 vccd1 vccd1 _4630__398/HI net398 sky130_fd_sc_hd__conb_1
XFILLER_0_9_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2290_ _0842_ _1067_ _0859_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3813_ net277 vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
XANTENNA_15 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2424__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_48 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3744_ net279 vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__inv_2
XANTENNA_59 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3675_ net241 vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2626_ _0828_ _1117_ _1132_ _1235_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a31o_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2557_ _1239_ _1241_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2488_ net706 net132 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\] vssd1
+ vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__a22o_1
X_4227_ clknet_leaf_47_wb_clk_i team_10_WB.instance_to_wrap.host_message_reg.next_state
+ _0216_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.Cstate
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ clknet_leaf_44_wb_clk_i net554 _0147_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3109_ team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked _0893_ net224 vssd1 vssd1
+ vccd1 vccd1 _1548_ sky130_fd_sc_hd__and3_4
X_4089_ clknet_leaf_8_wb_clk_i _0560_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2014__A3 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2486__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2238__B1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput24 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2260__A team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2961__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3460_ team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] net173 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[78\]
+ _0821_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2411_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__or4b_1
X_3391_ team_10_WB.instance_to_wrap.host_row2\[51\] net168 _1703_ team_10_WB.instance_to_wrap.host_row1\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2342_ _0820_ _0864_ _0842_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2273_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _0798_ _0801_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__o22a_1
X_4012_ clknet_leaf_32_wb_clk_i _0500_ net271 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2477__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2419__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2435__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4776_ net181 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1988_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] net148 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3727_ net241 vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2952__B2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3658_ net250 vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2609_ _0886_ _1274_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3589_ net284 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__inv_2
XANTENNA__2704__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1994__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2459__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _0994_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
XANTENNA__3120__A1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2960_ net125 _1482_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__nand2_2
XFILLER_0_130_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1911_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\] vssd1 vssd1 vccd1 vccd1
+ _0834_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2891_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] net1 _1227_ vssd1 vssd1 vccd1
+ vccd1 _1471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4630_ net398 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_71_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4561_ net372 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3512_ net235 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4492_ clknet_leaf_55_wb_clk_i _0017_ _0475_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3443_ team_10_WB.instance_to_wrap.host_row2\[53\] net168 net165 team_10_WB.instance_to_wrap.host_row2\[77\]
+ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3374_ _1747_ _1750_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2325_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1858_ vssd1 vssd1 vccd1 vccd1
+ _1101_ sky130_fd_sc_hd__or4b_1
XFILLER_0_97_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3025__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2256_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] net213 vssd1 vssd1 vccd1
+ vccd1 _1038_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2187_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net212 vssd1 vssd1 vccd1
+ vccd1 _0976_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3414__A2 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4759_ net180 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4562__373 vssd1 vssd1 vccd1 vccd1 _4562__373/HI net373 sky130_fd_sc_hd__conb_1
XFILLER_0_136_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3169__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1922__A_N net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2110_ team_10_WB.instance_to_wrap.dispFSM.guesses\[2\] net110 net134 net788 vssd1
+ vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__o22a_1
Xhold2 team_10_WB.instance_to_wrap.keypadFSMHost.strobe vssd1 vssd1 vccd1 vccd1 net554
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3090_ net199 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] net185 _1539_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[81\] sky130_fd_sc_hd__a31o_1
XFILLER_0_94_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2041_ team_10_WB.instance_to_wrap.dispFSM.guesses\[79\] net142 net108 net747 vssd1
+ vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3992_ clknet_leaf_44_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[29\]
+ _0060_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2943_ net736 net156 vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3809__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1958__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2874_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] _1459_ vssd1 vssd1 vccd1
+ vccd1 _1460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4613_ team_10_WB.instance_to_wrap.blue vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4544_ net355 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4475_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[32\]
+ _0458_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3426_ team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.dispFSM.guesses\[69\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3357_ team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] net168 net167 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2308_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] _1078_ _1083_
+ _1082_ _1079_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__o32a_1
XFILLER_0_77_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3288_ net741 _1671_ net228 vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__o21ai_1
X_2239_ _0796_ net208 _0799_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _1020_
+ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4546__357 vssd1 vssd1 vccd1 vccd1 _4546__357/HI net357 sky130_fd_sc_hd__conb_1
XFILLER_0_14_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3719__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold304_A team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input22_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2590_ net193 _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2_2
XFILLER_0_23_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4260_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[3\]
+ _0249_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3211_ net170 _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4191_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[53\]
+ _0180_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[53\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3142_ _1286_ _1554_ _1556_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__and3b_1
X_3073_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\]
+ net185 vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__mux2_1
X_2024_ _0904_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3975_ clknet_leaf_43_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[12\]
+ _0043_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2926_ net729 net154 net124 net676 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[31\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2857_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\] _1448_ vssd1 vssd1
+ vccd1 vccd1 _1450_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2788_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1397_ vssd1 vssd1 vccd1 vccd1
+ _1398_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_5_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold210 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\] vssd1 vssd1 vccd1
+ vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4527_ net338 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
Xhold221 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\] vssd1 vssd1 vccd1
+ vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] vssd1 vssd1 vccd1
+ vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\] vssd1 vssd1 vccd1
+ vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\] vssd1 vssd1 vccd1 vccd1
+ net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold265 team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] vssd1 vssd1 vccd1 vccd1
+ net817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\] vssd1 vssd1 vccd1
+ vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ clknet_leaf_46_wb_clk_i net720 _0441_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold287 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\] vssd1 vssd1 vccd1
+ vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold298 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] vssd1 vssd1 vccd1
+ vccd1 net850 sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ team_10_WB.instance_to_wrap.host_row1\[44\] _1693_ net171 team_10_WB.instance_to_wrap.host_row2\[84\]
+ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__a22o_1
X_4389_ clknet_leaf_4_wb_clk_i _0774_ _0372_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3069__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_105 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_116 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_127 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741__509 vssd1 vssd1 vccd1 vccd1 _4741__509/HI net509 sky130_fd_sc_hd__conb_1
XFILLER_0_113_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4635__403 vssd1 vssd1 vccd1 vccd1 _4635__403/HI net403 sky130_fd_sc_hd__conb_1
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3912__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3760_ net291 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2711_ net737 _1345_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3691_ net276 vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2642_ net215 _0952_ _1306_ _0951_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[1\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2573_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\] _1257_ vssd1 vssd1
+ vccd1 vccd1 _1258_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4312_ clknet_leaf_15_wb_clk_i _0702_ _0301_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4243_ clknet_leaf_48_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[7\]
+ _0232_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4174_ clknet_leaf_46_wb_clk_i _0643_ _0163_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3125_ _0824_ _1861_ _1555_ _1291_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3033__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3056_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] _1522_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\] sky130_fd_sc_hd__mux2_2
XFILLER_0_78_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2007_ net216 net217 vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2274__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3471__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3958_ clknet_leaf_47_wb_clk_i _0009_ _0026_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2909_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\] net151 net122 net833
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[14\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3889_ net261 vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3453__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3812_ net290 vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__inv_2
XANTENNA_16 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3743_ net279 vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3674_ net269 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2625_ _0010_ _0007_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[1\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput101 net181 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2556_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] _1243_ _1245_
+ _1242_ _1239_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2487_ net616 net129 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1
+ vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4226_ clknet_leaf_10_wb_clk_i net534 _0215_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[101\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4157_ clknet_leaf_45_wb_clk_i net556 _0146_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3108_ net82 net40 net42 vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__and3b_1
XFILLER_0_39_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4088_ clknet_leaf_9_wb_clk_i _0559_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3039_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\]
+ net185 vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3444__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2798__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2014__A4 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4747__515 vssd1 vssd1 vccd1 vccd1 _4747__515/HI net515 sky130_fd_sc_hd__conb_1
XFILLER_0_92_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2806__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2238__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1997__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput14 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput36 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2260__B _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2410_ team_10_WB.instance_to_wrap.clock_div.count\[2\] team_10_WB.instance_to_wrap.clock_div.count\[4\]
+ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or3_1
X_3390_ _1763_ _1765_ _1766_ net302 vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__o31a_1
XFILLER_0_122_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2341_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _1112_ _1115_ vssd1 vssd1
+ vccd1 vccd1 _1117_ sky130_fd_sc_hd__and3b_1
XFILLER_0_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2272_ _0792_ net211 _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1
+ vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__a22o_1
XANTENNA__3091__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4011_ clknet_leaf_32_wb_clk_i _0499_ net271 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_75_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3426__A0 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2435__B _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1988__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4775_ net182 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
X_1987_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net147 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3726_ net252 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout122_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3657_ net264 vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2608_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\] _1275_ _1284_ _1289_
+ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3588_ net269 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__inv_2
XANTENNA__2165__A0 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2539_ team_10_WB.instance_to_wrap.host_col\[3\] _0852_ _1179_ vssd1 vssd1 vccd1
+ vccd1 _0487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3282__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4209_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[71\]
+ _0198_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[71\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1979__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2459__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 net182 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
XANTENNA__3920__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 _1222_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4058__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3408__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2255__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1910_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\] vssd1 vssd1 vccd1 vccd1
+ _0833_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2890_ net191 _1470_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_31_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4560_ net371 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3511_ net235 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4491_ clknet_leaf_47_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_state _0474_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.Cstate sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3442_ _1800_ _1813_ _1815_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3373_ team_10_WB.instance_to_wrap.host_row1\[66\] _1703_ net178 team_10_WB.instance_to_wrap.host_row2\[58\]
+ _1748_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2324_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2255_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net211 vssd1 vssd1 vccd1
+ vccd1 _1037_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2186_ _0822_ _0952_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3041__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4758_ net180 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2925__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3709_ net232 vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4689_ net457 vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_2
XFILLER_0_120_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2138__A0 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3341__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold3 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge vssd1 vssd1 vccd1 vccd1
+ net555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ team_10_WB.instance_to_wrap.dispFSM.guesses\[72\] net113 net137 team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3991_ clknet_leaf_44_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[28\]
+ _0059_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2942_ net208 net154 net124 net684 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[47\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2873_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net221 vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__or3b_1
XANTENNA__3097__A team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4612_ net386 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_2_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2907__A2 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4543_ net354 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4474_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[31\]
+ _0457_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3425_ team_10_WB.instance_to_wrap.host_row1\[45\] net302 _1693_ vssd1 vssd1 vccd1
+ vccd1 _1800_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3036__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2032__B1_N net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3332__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3356_ team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] net165 _1732_ _1734_ vssd1
+ vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2307_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__inv_2
X_3287_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\] _1671_ vssd1 vssd1 vccd1
+ vccd1 _1672_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout287_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2238_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _0804_ _0800_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ team_10_WB.instance_to_wrap.correct\[0\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4003__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3210_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ _1621_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4190_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[52\]
+ _0179_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[52\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3141_ _1563_ _1570_ _0905_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3072_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] _1530_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[72\] sky130_fd_sc_hd__mux2_1
X_2023_ _0893_ _0895_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3974_ clknet_leaf_42_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[11\]
+ _0042_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2925_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\] net151 net122 net795
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[30\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__2443__B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2053__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2856_ _1448_ _1449_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2787_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__and4b_1
XFILLER_0_108_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3555__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold200 team_10_WB.instance_to_wrap.dispFSM.guesses\[67\] vssd1 vssd1 vccd1 vccd1
+ net752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 team_10_WB.instance_to_wrap.dispFSM.guesses\[77\] vssd1 vssd1 vccd1 vccd1
+ net763 sky130_fd_sc_hd__dlygate4sd3_1
X_4526_ net337 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout202_A team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold222 team_10_WB.instance_to_wrap.dispFSM.guesses\[44\] vssd1 vssd1 vccd1 vccd1
+ net774 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold233 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\] vssd1 vssd1 vccd1
+ vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\] vssd1 vssd1 vccd1
+ vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\] vssd1 vssd1 vccd1
+ vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4457_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[14\]
+ _0440_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] vssd1 vssd1 vccd1 vccd1
+ net818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold277 team_10_WB.instance_to_wrap.clock_div.count\[15\] vssd1 vssd1 vccd1 vccd1
+ net829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 team_10_WB.instance_to_wrap.dispFSM.guesses\[12\] vssd1 vssd1 vccd1 vccd1
+ net840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 team_10_WB.instance_to_wrap.clock_div.count\[20\] vssd1 vssd1 vccd1 vccd1
+ net851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3408_ team_10_WB.instance_to_wrap.host_row1\[52\] _1699_ net165 team_10_WB.instance_to_wrap.host_row2\[76\]
+ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4388_ clknet_leaf_23_wb_clk_i _0773_ _0371_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_input7_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3339_ _1687_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__nor2_4
X_4513__324 vssd1 vssd1 vccd1 vccd1 _4513__324/HI net324 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_106 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_117 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_139 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4674__442 vssd1 vssd1 vccd1 vccd1 _4674__442/HI net442 sky130_fd_sc_hd__conb_1
XFILLER_0_20_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2504__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4715__483 vssd1 vssd1 vccd1 vccd1 _4715__483/HI net483 sky130_fd_sc_hd__conb_1
XFILLER_0_21_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2809__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4181__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2710_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3690_ net231 vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2641_ _0945_ _1305_ _0936_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2572_ net216 net224 vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4311_ clknet_leaf_14_wb_clk_i _0701_ _0300_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4242_ clknet_leaf_48_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[6\]
+ _0231_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4173_ clknet_leaf_46_wb_clk_i _0642_ _0162_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_138_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3124_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3055_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\]
+ net185 vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2006_ net216 net217 vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2274__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout152_A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ clknet_leaf_45_wb_clk_i _0008_ _0025_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2908_ net694 net154 net124 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[13\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3888_ net261 vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4658__426 vssd1 vssd1 vccd1 vccd1 _4658__426/HI net426 sky130_fd_sc_hd__conb_1
X_2839_ _0518_ _1439_ _1436_ _1411_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4509_ net320 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4091__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3089__B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3811_ net273 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_17 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_28 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3742_ net291 vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3673_ net264 vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2624_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] _1074_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_3_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2555_ _1246_ _1239_ _1244_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__and3b_1
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2486_ net678 net129 net125 team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\] _1190_
+ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__a221o_1
X_4225_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[87\]
+ _0214_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[87\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4156_ clknet_leaf_38_wb_clk_i _0627_ net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3107_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1395_ _1547_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.lcd_en sky130_fd_sc_hd__nor3_1
XFILLER_0_78_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4087_ clknet_leaf_8_wb_clk_i _0558_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3038_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] _1513_ net200 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[55\] sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2247__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2955__B1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4519__330 vssd1 vssd1 vccd1 vccd1 _4519__330/HI net330 sky130_fd_sc_hd__conb_1
XFILLER_0_44_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4574__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1997__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4606__380 vssd1 vssd1 vccd1 vccd1 _4606__380/HI net380 sky130_fd_sc_hd__conb_1
XFILLER_0_68_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput15 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput26 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput37 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3371__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2340_ _1112_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2271_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] _0803_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ _1048_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__o221a_1
XANTENNA__2269__A team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4010_ clknet_leaf_33_wb_clk_i _0498_ net271 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_79_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2477__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4774_ net529 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1986_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] _0874_ _0882_ net156 vssd1
+ vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2937__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3725_ net253 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3039__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3656_ net271 vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2607_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1288_ _1270_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3587_ net269 vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3362__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2538_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0840_ _1235_ vssd1 vssd1
+ vccd1 vccd1 _0504_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2469_ net808 net130 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\]
+ _1208_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__a221o_1
X_4208_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[70\]
+ _0197_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[70\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4139_ clknet_leaf_3_wb_clk_i _0610_ _0138_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1979__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2928__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3353__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout170 _1612_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
XANTENNA__2459__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout181 net182 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xfanout192 _0991_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2919__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3510_ net235 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4490_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[47\]
+ _0473_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3441_ net178 _1802_ _1809_ _1701_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3344__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3372_ team_10_WB.instance_to_wrap.host_row2\[50\] net168 net177 team_10_WB.instance_to_wrap.host_row2\[66\]
+ _1749_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2323_ _1097_ _1098_ _0868_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__a21oi_1
X_2254_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net211 vssd1 vssd1 vccd1
+ vccd1 _1036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2185_ net133 _0972_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4757_ net525 vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_2
X_1969_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] net147 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\]
+ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2386__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3708_ net232 vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4688_ net456 vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_2
XFILLER_0_4_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3639_ net285 vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3102__A3 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3326__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge vssd1 vssd1 vccd1 vccd1
+ net556 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2301__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2266__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ clknet_leaf_45_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[27\]
+ _0058_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2941_ net209 net151 net122 net772 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[46\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2872_ _1222_ _1458_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[0\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4611_ net385 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_13_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3014__C1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4542_ net353 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4473_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[30\]
+ _0456_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4691__459 vssd1 vssd1 vccd1 vccd1 _4691__459/HI net459 sky130_fd_sc_hd__conb_1
XFILLER_0_110_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3424_ team_10_WB.instance_to_wrap.host_row1\[77\] net301 _1708_ vssd1 vssd1 vccd1
+ vccd1 _1799_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4619__390 vssd1 vssd1 vccd1 vccd1 _4619__390/HI net390 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3355_ team_10_WB.instance_to_wrap.dispFSM.guesses\[65\] _1719_ _1733_ net229 vssd1
+ vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__a211o_1
XANTENNA__3841__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2306_ _0841_ _1073_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__or2_2
X_3286_ net294 _1670_ _1671_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__nor3_1
X_2237_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _0799_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\]
+ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__a221o_1
XANTENNA__3052__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2168_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2099_ net696 net143 net107 net698 vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4626__394 vssd1 vssd1 vccd1 vccd1 _4626__394/HI net394 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3020__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4048__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2522__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3140_ _0889_ _0894_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3071_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\]
+ net185 vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2022_ _0892_ _0896_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2038__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3973_ clknet_leaf_42_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[10\]
+ _0041_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2924_ net672 net154 net124 net657 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[29\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2855_ net744 _1447_ net174 vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2786_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1 _1396_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_48_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4525_ net336 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
Xhold201 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\] vssd1 vssd1 vccd1 vccd1
+ net753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2210__B1 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\] vssd1 vssd1 vccd1 vccd1
+ net764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3047__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold223 team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] vssd1 vssd1 vccd1 vccd1
+ net775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] vssd1 vssd1 vccd1 vccd1
+ net786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold245 team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] vssd1 vssd1 vccd1 vccd1
+ net797 sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ clknet_leaf_26_wb_clk_i net695 _0439_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold256 team_10_WB.instance_to_wrap.host_row1\[58\] vssd1 vssd1 vccd1 vccd1 net808
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] vssd1 vssd1 vccd1
+ vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold278 team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\] vssd1 vssd1 vccd1 vccd1
+ net830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3407_ net67 net175 _1783_ net228 vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold289 team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] vssd1 vssd1 vccd1 vccd1
+ net841 sky130_fd_sc_hd__dlygate4sd3_1
X_4387_ clknet_leaf_22_wb_clk_i _0772_ _0370_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_102_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3338_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net206 _1707_ vssd1 vssd1
+ vccd1 vccd1 _1718_ sky130_fd_sc_hd__or3_2
X_4552__363 vssd1 vssd1 vccd1 vccd1 _4552__363/HI net363 sky130_fd_sc_hd__conb_1
XFILLER_0_119_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3269_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\]
+ _1657_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_107 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_118 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_129 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2268__B1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2825__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3480__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2440__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2640_ _0926_ net185 vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__nand2_1
XANTENNA__2991__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4495__306 vssd1 vssd1 vccd1 vccd1 _4495__306/HI net306 sky130_fd_sc_hd__conb_1
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2571_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] _0898_ vssd1 vssd1
+ vccd1 vccd1 _1256_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4310_ clknet_leaf_30_wb_clk_i _0700_ _0299_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[33\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4241_ clknet_leaf_48_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[5\]
+ _0230_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] sky130_fd_sc_hd__dfrtp_1
X_4536__347 vssd1 vssd1 vccd1 vccd1 _4536__347/HI net347 sky130_fd_sc_hd__conb_1
XFILLER_0_103_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4172_ clknet_leaf_46_wb_clk_i _0641_ _0161_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3123_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] _1288_ _1553_ _0825_
+ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3054_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] _1521_ net200 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[63\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ net217 net219 net220 vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__or3_2
XFILLER_0_52_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3471__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2454__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3956_ clknet_leaf_45_wb_clk_i _0007_ _0024_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout145_A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2907_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\] net152 net123 net766
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[12\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3887_ net261 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4697__465 vssd1 vssd1 vccd1 vccd1 _4697__465/HI net465 sky130_fd_sc_hd__conb_1
X_2838_ _1407_ _0515_ _1426_ _1409_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__o31a_1
XFILLER_0_85_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2769_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[25\]
+ team_10_WB.instance_to_wrap.clock_div.count\[24\] _1380_ vssd1 vssd1 vccd1 vccd1
+ _1384_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4508_ net319 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_112_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4439_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[36\]
+ _0422_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3462__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3150__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3810_ net290 vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3741_ net278 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2964__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3672_ net274 vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2623_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1074_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2554_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] _1241_ vssd1 vssd1 vccd1
+ vccd1 _1246_ sky130_fd_sc_hd__and4_1
XFILLER_0_122_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2485_ net726 net132 _1187_ _1215_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4224_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[86\]
+ _0213_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[86\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4155_ clknet_leaf_44_wb_clk_i _0626_ _0145_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3106_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ _1546_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] vssd1 vssd1 vccd1 vccd1
+ _1547_ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ clknet_leaf_8_wb_clk_i _0557_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3037_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3444__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3939_ net270 vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4786__533 vssd1 vssd1 vccd1 vccd1 _4786__533/HI net533 sky130_fd_sc_hd__conb_1
XFILLER_0_22_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1997__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput16 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3934__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2270_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net209 vssd1 vssd1 vccd1
+ vccd1 _1052_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2269__B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1988__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4773_ net180 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] net145 vssd1 vssd1 vccd1
+ vccd1 _0882_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2937__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3724_ net253 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3655_ net258 vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2606_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] _1287_ vssd1 vssd1
+ vccd1 vccd1 _1288_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3586_ net287 vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4081__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2537_ _0871_ _1073_ _1088_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__nand3_1
XANTENNA__3055__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2468_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] net195 vssd1 vssd1
+ vccd1 vccd1 _1208_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3114__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4207_ clknet_leaf_32_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[69\]
+ _0196_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[69\] sky130_fd_sc_hd__dfrtp_1
X_2399_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[6\]
+ team_10_WB.instance_to_wrap.clock_div.count\[5\] vssd1 vssd1 vccd1 vccd1 _1162_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_39_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4138_ clknet_leaf_24_wb_clk_i _0609_ _0137_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4069_ clknet_leaf_36_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[0\]
+ _0089_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3417__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1979__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3050__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4753__521 vssd1 vssd1 vccd1 vccd1 _4753__521/HI net521 sky130_fd_sc_hd__conb_1
XFILLER_0_104_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input38_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4585__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 net161 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_2
Xfanout171 _1701_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_4
Xfanout182 net101 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_2
Xfanout193 _0885_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3408__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3929__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3440_ _1707_ _1804_ _1814_ _1717_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3371_ team_10_WB.instance_to_wrap.host_row2\[82\] net171 _1708_ team_10_WB.instance_to_wrap.host_row1\[74\]
+ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2322_ _0844_ _0851_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2253_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] net210 vssd1 vssd1 vccd1
+ vccd1 _1035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2184_ _0919_ _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4756_ net524 vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_2
XFILLER_0_16_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1968_ net743 net148 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] vssd1
+ vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4737__505 vssd1 vssd1 vccd1 vccd1 _4737__505/HI net505 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3707_ net232 vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__inv_2
X_4687_ net455 vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_2
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1899_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _0823_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3638_ net285 vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3569_ net244 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold5 team_10_WB.instance_to_wrap.clock_div.count\[29\] vssd1 vssd1 vccd1 vccd1 net557
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2940_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] net155 _1472_ net680 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[45\] sky130_fd_sc_hd__a22o_1
XFILLER_0_85_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2871_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] _1457_ vssd1 vssd1 vccd1
+ vccd1 _1458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4610_ net384 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4541_ net352 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_53_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4472_ clknet_leaf_33_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[29\]
+ _0455_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3423_ net68 net176 _1798_ net227 vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4591__550 vssd1 vssd1 vccd1 vccd1 net550 _4591__550/LO sky130_fd_sc_hd__conb_1
XFILLER_0_81_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3354_ team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] net171 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2305_ _0841_ _0860_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_1
X_3285_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\]
+ _1666_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2236_ _0796_ net208 net211 _0797_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__a22o_1
XANTENNA__3096__A3 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2167_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2098_ team_10_WB.instance_to_wrap.dispFSM.guesses\[14\] net114 net137 net841 vssd1
+ vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4739_ net507 vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_2
XFILLER_0_90_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3244__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output69_A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3070_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _1529_ net201 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[71\] sky130_fd_sc_hd__mux2_1
X_2021_ _0892_ _0894_ net225 vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__or3b_2
XFILLER_0_82_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3972_ clknet_leaf_43_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[9\]
+ _0040_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2923_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\] net152 net123 net815
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[28\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2854_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ _1444_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2785_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\]
+ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4524_ net335 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
Xhold202 team_10_WB.instance_to_wrap.dispFSM.guesses\[19\] vssd1 vssd1 vccd1 vccd1
+ net754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold213 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] vssd1 vssd1 vccd1
+ vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\] vssd1 vssd1 vccd1
+ vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 team_10_WB.instance_to_wrap.gamelogic.rights\[1\] vssd1 vssd1 vccd1 vccd1
+ net798 sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[12\]
+ _0438_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold257 team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] vssd1 vssd1 vccd1 vccd1
+ net809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold279 team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] vssd1 vssd1 vccd1 vccd1
+ net831 sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ net229 _1774_ _1782_ _1767_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__a211o_1
X_4386_ clknet_leaf_47_wb_clk_i _0771_ _0369_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3337_ _1694_ _1714_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout292_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3063__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3268_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ net739 vssd1 vssd1
+ vccd1 vccd1 _1659_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2187__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2219_ net28 net29 vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__nand2_1
X_3199_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] _1392_ vssd1 vssd1 vccd1
+ vccd1 _1617_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3474__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_108 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_119 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2201__A1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3762__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input20_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2268__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2955__A2_N _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2570_ net220 net224 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] vssd1
+ vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3672__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4240_ clknet_leaf_50_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[4\]
+ _0229_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4171_ clknet_leaf_46_wb_clk_i _0640_ _0160_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_120_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3122_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\] _1552_ _0824_ vssd1
+ vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3053_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__mux2_1
XANTENNA__2259__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3456__B1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2004_ net300 net3 vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3955_ clknet_leaf_45_wb_clk_i _0006_ _0023_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2906_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\] net151 net122 net767
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[11\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3886_ net260 vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2837_ _1407_ _1436_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3058__S net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2768_ team_10_WB.instance_to_wrap.clock_div.count\[24\] _1382_ net826 vssd1 vssd1
+ vccd1 vccd1 _1383_ sky130_fd_sc_hd__a21oi_1
X_4507_ net318 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_41_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2699_ _0807_ team_10_WB.instance_to_wrap.message_reg.state\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ _1343_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _1344_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4438_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[35\]
+ _0421_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4369_ clknet_leaf_20_wb_clk_i _0754_ _0352_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_22_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3447__B1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2645__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3667__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_19 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3740_ net292 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4503__314 vssd1 vssd1 vccd1 vccd1 _4503__314/HI net314 sky130_fd_sc_hd__conb_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3671_ net256 vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2622_ _1116_ _1235_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_23_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2553_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2484_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\] _0991_ vssd1 vssd1 vccd1
+ vccd1 _1215_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4223_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[85\]
+ _0212_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[85\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4154_ clknet_leaf_9_wb_clk_i _0625_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3105_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1396_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_78_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4085_ clknet_leaf_8_wb_clk_i _0556_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3036_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _1512_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[54\] sky130_fd_sc_hd__mux2_1
XFILLER_0_78_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2465__B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2101__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4664__432 vssd1 vssd1 vccd1 vccd1 _4664__432/HI net432 sky130_fd_sc_hd__conb_1
XFILLER_0_17_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout255_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4705__473 vssd1 vssd1 vccd1 vccd1 _4705__473/HI net473 sky130_fd_sc_hd__conb_1
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3938_ net253 vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3869_ net283 vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2891__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3487__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput17 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput28 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput39 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3426__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3371__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4648__416 vssd1 vssd1 vccd1 vccd1 _4648__416/HI net416 sky130_fd_sc_hd__conb_1
XFILLER_0_75_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4772_ net180 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1984_ net761 net147 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1
+ vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2937__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3723_ net253 vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3654_ net258 vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2605_ _0888_ _1279_ _0900_ _0899_ _0895_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_24_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3585_ net284 vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3362__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2536_ net580 team_10_WB.instance_to_wrap.buffer.temp_guess\[0\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2467_ net612 net128 _1207_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4206_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\]
+ _0195_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[68\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2398_ team_10_WB.instance_to_wrap.clock_div.count\[8\] team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] vssd1 vssd1 vccd1 vccd1 _1161_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4137_ clknet_leaf_20_wb_clk_i _0608_ _0136_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3071__S net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4068_ clknet_leaf_51_wb_clk_i _0550_ _0088_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_78_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3019_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] net189 vssd1 vssd1 vccd1
+ vccd1 _1504_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3353__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2561__B1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout150 net152 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
Xfanout172 _1696_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout183 _0995_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xfanout194 _0855_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2092__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3370_ team_10_WB.instance_to_wrap.host_row1\[42\] _1693_ net172 team_10_WB.instance_to_wrap.host_row2\[42\]
+ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__a22o_1
XANTENNA__3344__A2 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2321_ _0819_ _0849_ _0851_ _0867_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__or4_1
XFILLER_0_85_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2252_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] _1033_ _1025_ _1027_
+ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_109_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2183_ _0923_ _0947_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4509__320 vssd1 vssd1 vccd1 vccd1 _4509__320/HI net320 sky130_fd_sc_hd__conb_1
XFILLER_0_8_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4755_ net523 vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1967_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] net147 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3706_ net232 vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout120_A _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4686_ net454 vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_2
XFILLER_0_31_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1898_ net215 vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3637_ net264 vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3568_ net244 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2519_ net619 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] vssd1 vssd1
+ vccd1 vccd1 _0526_ sky130_fd_sc_hd__a22o_1
X_3499_ net235 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3326__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4596__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold6 team_10_WB.instance_to_wrap.gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 net558
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2870_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net221 vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4540_ net351 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4471_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[28\]
+ _0454_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3422_ net229 _1788_ _1794_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3353_ team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] net178 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[9\]
+ _1731_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2304_ _0868_ _1080_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__o21a_1
X_3284_ net820 _1668_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2235_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _0800_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2166_ _0936_ _0939_ _0954_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2097_ net687 net142 net108 net693 vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2461__C1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3005__B2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2999_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\] net159 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[32\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4738_ net506 vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_2
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4669_ net437 vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_2
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4094__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3434__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2020_ _0899_ _0902_ _0901_ _0896_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_136_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3971_ clknet_leaf_43_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[8\]
+ _0039_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2922_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\] net150 net121 net807
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[27\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2853_ _1447_ net174 _1446_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[4\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_45_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2784_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4523_ net334 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold203 team_10_WB.instance_to_wrap.dispFSM.guesses\[79\] vssd1 vssd1 vccd1 vccd1
+ net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\] vssd1 vssd1 vccd1
+ vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold225 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\] vssd1 vssd1 vccd1
+ vccd1 net777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold236 team_10_WB.instance_to_wrap.dispFSM.guesses\[10\] vssd1 vssd1 vccd1 vccd1
+ net788 sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[11\]
+ _0437_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold247 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\] vssd1 vssd1 vccd1 vccd1
+ net799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] vssd1 vssd1 vccd1
+ vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] vssd1 vssd1 vccd1 vccd1
+ net821 sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\] _1690_ net173 _1775_
+ _1781_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__a221o_1
X_4385_ clknet_leaf_3_wb_clk_i _0770_ _0368_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] net165 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[72\]
+ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__a22o_1
XANTENNA__2468__B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3267_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ _1658_ vssd1 vssd1
+ vccd1 vccd1 _0561_ sky130_fd_sc_hd__o21a_1
X_2218_ net25 net24 net27 net26 vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3198_ _1393_ _1611_ _1616_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_109 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2149_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] _0943_ vssd1 vssd1 vccd1
+ vccd1 _0944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3465__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2268__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input13_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4681__449 vssd1 vssd1 vccd1 vccd1 _4681__449/HI net449 sky130_fd_sc_hd__conb_1
XFILLER_0_129_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2440__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2569__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4170_ clknet_leaf_46_wb_clk_i _0639_ _0159_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_3121_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] _1860_ vssd1 vssd1
+ vccd1 vccd1 _1552_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3052_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] _1520_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[62\] sky130_fd_sc_hd__mux2_1
XFILLER_0_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2259__A2 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3977__CLK clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1920__B net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2003_ team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3954_ clknet_leaf_47_wb_clk_i _0005_ _0022_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2905_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\] net151 net122 net769
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[10\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3885_ net283 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2836_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2767_ net715 _1382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[24\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4506_ net317 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_48_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3392__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2698_ team_10_WB.instance_to_wrap.message_reg.msg\[0\] team_10_WB.instance_to_wrap.message_reg.msg\[1\]
+ team_10_WB.instance_to_wrap.message_reg.msg\[2\] team_10_WB.instance_to_wrap.message_reg.msg\[3\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4437_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[34\]
+ _0420_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3074__S net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4368_ clknet_leaf_46_wb_clk_i _0753_ _0351_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input5_A gpio_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3319_ _1688_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__and2_4
X_4299_ clknet_leaf_13_wb_clk_i _0689_ _0288_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_119_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2587__A1_N net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2489__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3438__A1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3438__B2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2949__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4542__353 vssd1 vssd1 vccd1 vccd1 _4542__353/HI net353 sky130_fd_sc_hd__conb_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3670_ net254 vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2621_ _0006_ _0009_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_109_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3683__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2552_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] _1243_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_23_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2483_ net641 net131 _1185_ _1214_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4222_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[84\]
+ _0211_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[84\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4153_ clknet_leaf_12_wb_clk_i _0624_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3104_ team_10_WB.EN_VAL_REG net181 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__or2_1
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4084_ clknet_leaf_8_wb_clk_i _0555_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3429__A1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3035_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout150_A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3937_ net253 vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__inv_2
X_4779__531 vssd1 vssd1 vccd1 vccd1 _4779__531/HI net531 sky130_fd_sc_hd__conb_1
XFILLER_0_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3069__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3868_ net287 vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2819_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3799_ net279 vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2701__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_55_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4526__337 vssd1 vssd1 vccd1 vccd1 _4526__337/HI net337 sky130_fd_sc_hd__conb_1
XFILLER_0_49_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4687__455 vssd1 vssd1 vccd1 vccd1 _4687__455/HI net455 sky130_fd_sc_hd__conb_1
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4728__496 vssd1 vssd1 vccd1 vccd1 _4728__496/HI net496 sky130_fd_sc_hd__conb_1
XFILLER_0_75_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4771_ net528 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
X_1983_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] _0874_ _0881_ net156 vssd1
+ vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3722_ net252 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3653_ net287 vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2604_ _1268_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\] _1265_ vssd1
+ vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__or3b_2
XFILLER_0_70_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3584_ net264 vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2535_ net582 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2570__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2466_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] net196 _1187_
+ _1206_ net131 vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4205_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[67\]
+ _0194_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[67\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2397_ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ team_10_WB.instance_to_wrap.clock_div.count\[9\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__or4bb_1
XANTENNA_fanout198_A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4136_ clknet_leaf_27_wb_clk_i _0607_ _0135_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2476__B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4067_ clknet_leaf_50_wb_clk_i _0549_ _0087_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3018_ net195 _1503_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[45\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_78_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout140 _0914_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_4
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout173 _1696_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_2
Xfanout184 _0995_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
Xfanout195 _0826_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2077__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4006__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2001__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2320_ _1094_ _1095_ _0869_ _1092_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2251_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0798_ _0800_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\]
+ _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2182_ net215 net214 team_10_WB.instance_to_wrap.gamelogic.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _0971_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2068__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4754_ net522 vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1966_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0874_ _0878_ net158 vssd1
+ vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ net233 vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4685_ net453 vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_2
XFILLER_0_16_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1897_ net299 vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3636_ net249 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3567_ net276 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3871__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2518_ _0807_ _0808_ net142 vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__and3_2
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3498_ net276 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2449_ net630 net132 _1191_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3082__S net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4119_ clknet_leaf_5_wb_clk_i _0590_ _0118_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3008__C1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input43_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold7 team_10_WB.instance_to_wrap.host_row1\[101\] vssd1 vssd1 vccd1 vccd1 net559
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3014__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4470_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[27\]
+ _0453_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3421_ net177 _1795_ _1796_ net173 _1781_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__a221o_1
XANTENNA__4787__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2525__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3352_ team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] net172 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[73\]
+ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2303_ net222 net223 _0869_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__or3_1
X_3283_ net625 _1666_ _1669_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2234_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] _0805_ vssd1 vssd1 vccd1
+ vccd1 _1016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2165_ _0942_ _0955_ net872 vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2096_ team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] net113 net137 net794 vssd1
+ vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__o22a_1
X_4743__511 vssd1 vssd1 vccd1 vccd1 _4743__511/HI net511 sky130_fd_sc_hd__conb_1
XFILLER_0_49_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3005__A2 net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2998_ net125 _1496_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__nand2_2
XFILLER_0_133_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4737_ net505 vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1949_ _0841_ _0871_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3077__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4668_ net436 vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_2
XFILLER_0_102_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3619_ net244 vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4599_ net197 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3477__C1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2945__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1963__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3468__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3483__A2 _1853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3970_ clknet_leaf_43_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[7\]
+ _0038_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2921_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\] net152 net123 net771
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[26\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3686__A net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2590__A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2852_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\]
+ _1442_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2783_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4522_ net333 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_108_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold204 _0746_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold215 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\] vssd1 vssd1 vccd1
+ vccd1 net767 sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[10\]
+ _0436_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\]
+ sky130_fd_sc_hd__dfstp_1
Xhold226 team_10_WB.instance_to_wrap.dispFSM.guesses\[66\] vssd1 vssd1 vccd1 vccd1
+ net778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\] vssd1 vssd1 vccd1 vccd1
+ net789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold248 team_10_WB.instance_to_wrap.dispFSM.guesses\[64\] vssd1 vssd1 vccd1 vccd1
+ net800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold259 team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] vssd1 vssd1 vccd1 vccd1
+ net811 sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _1777_ _1780_ net175 vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4384_ clknet_leaf_46_wb_clk_i _0769_ _0367_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3335_ _1687_ _1714_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ net293 vssd1 vssd1
+ vccd1 vccd1 _1658_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2217_ net15 net17 net18 net16 vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout180_A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3197_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1616_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3474__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2148_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nand2_1
XANTENNA__2484__B _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2079_ team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] net109 net134 net867 vssd1
+ vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2704__S net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1960__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4061__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2976__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output74_A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3153__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3120_ net193 _1550_ _1290_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3051_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3456__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2002_ team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3953_ clknet_3_1_0_wb_clk_i _0016_ net268 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2904_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\] net149 net120 net839
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[9\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3884_ net286 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2835_ _1415_ _1426_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2766_ _1381_ _1382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[23\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4505_ net316 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2697_ _1341_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\] vssd1 vssd1
+ vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4436_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[33\]
+ _0419_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_112_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4367_ clknet_leaf_20_wb_clk_i _0752_ _0350_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3318_ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__inv_2
X_4298_ clknet_leaf_27_wb_clk_i net697 _0287_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3249_ _1610_ _1647_ net294 vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2495__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3447__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3383__A1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3383__B2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2949__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2620_ _0840_ _0860_ _1295_ _1085_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2551_ _1239_ _1242_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_45_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2482_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] net184 vssd1 vssd1 vccd1
+ vccd1 _1214_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4221_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[83\]
+ _0210_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[83\] sky130_fd_sc_hd__dfrtp_1
X_4152_ clknet_leaf_12_wb_clk_i _0623_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_128_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3103_ net158 _1302_ net195 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_state
+ sky130_fd_sc_hd__mux2_1
X_4083_ clknet_leaf_8_wb_clk_i _0554_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3429__A2 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3034_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _1511_ net200 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[53\] sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3936_ net256 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3867_ net282 vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2818_ _1410_ _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3798_ net291 vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2749_ net852 _1370_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3085__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3117__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout300 net6 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
X_4419_ clknet_leaf_24_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[16\]
+ _0402_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold188_A team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3053__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_4
XFILLER_0_18_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1982_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] net145 vssd1 vssd1 vccd1
+ vccd1 _0881_ sky130_fd_sc_hd__or2_1
X_4770_ net180 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ net234 vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3652_ net248 vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2603_ _0016_ _0013_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[1\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3583_ net282 vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2534_ net568 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2465_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] net192 vssd1 vssd1 vccd1
+ vccd1 _1206_ sky130_fd_sc_hd__or2_1
X_4204_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[66\]
+ _0193_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[66\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2396_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0854_ _1158_ net656 vssd1
+ vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__a22o_1
X_4135_ clknet_leaf_11_wb_clk_i _0606_ _0134_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ clknet_leaf_51_wb_clk_i _0548_ _0086_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3017_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout260_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3035__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3919_ net242 vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2013__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout130 _1183_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout141 net143 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_2
Xfanout163 net164 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout174 _1440_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_2
Xfanout185 net187 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout196 _0826_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3019__A team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2001__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654__422 vssd1 vssd1 vccd1 vccd1 _4654__422/HI net422 sky130_fd_sc_hd__conb_1
XFILLER_0_122_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2250_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _0804_ _1029_ _1031_ vssd1
+ vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2181_ _0970_ team_10_WB.instance_to_wrap.correct\[0\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3689__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3017__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4753_ net521 vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_2
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1965_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] net144 vssd1 vssd1 vccd1
+ vccd1 _0878_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3704_ net232 vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4684_ net452 vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1896_ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3635_ net249 vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3566_ net276 vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2517_ team_10_WB.instance_to_wrap.message_reg.state\[1\] net142 _0808_ vssd1 vssd1
+ vccd1 vccd1 _1231_ sky130_fd_sc_hd__o21ai_4
X_3497_ net276 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2448_ net653 net131 _1187_ _1197_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2379_ _1099_ _1151_ _1135_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4118_ clknet_leaf_15_wb_clk_i _0589_ _0117_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4049_ clknet_leaf_7_wb_clk_i _0534_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4638__406 vssd1 vssd1 vccd1 vccd1 _4638__406/HI net406 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input36_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1 net560
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3247__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3021__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2470__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2470__B2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3420_ team_10_WB.instance_to_wrap.host_row2\[44\] team_10_WB.instance_to_wrap.dispFSM.guesses\[20\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3351_ net64 net175 _1730_ net228 vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2302_ _0844_ _0847_ _0853_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3282_ net294 _1668_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__nor2_1
X_2233_ _0797_ net211 _0804_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _1014_
+ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2164_ _0942_ _0943_ _0957_ _0955_ net830 vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2095_ team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] net109 net135 net712 vssd1
+ vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2461__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2997_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] _1494_ _1495_ vssd1
+ vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4736_ net504 vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_2
XFILLER_0_133_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1948_ _0865_ _0870_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nand2b_2
XANTENNA__3410__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4667_ net435 vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_2
X_1879_ net213 vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3618_ net244 vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4598_ net197 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3549_ net277 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3477__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2945__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2920_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\] net149 net120 net813
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[25\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2851_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] _1444_ vssd1 vssd1
+ vccd1 vccd1 _1446_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2782_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1392_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4521_ net332 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold205 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\] vssd1 vssd1 vccd1
+ vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold216 team_10_WB.instance_to_wrap.message_reg.state\[0\] vssd1 vssd1 vccd1 vccd1
+ net768 sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ clknet_leaf_47_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[9\]
+ _0435_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_83_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold227 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\] vssd1 vssd1 vccd1
+ vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold238 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\] vssd1 vssd1 vccd1
+ vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 team_10_WB.instance_to_wrap.dispFSM.guesses\[68\] vssd1 vssd1 vccd1 vccd1
+ net801 sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _1685_ _1720_ _1778_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4383_ clknet_leaf_1_wb_clk_i _0768_ _0366_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3334_ _1707_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net206 vssd1 vssd1
+ vccd1 vccd1 _1714_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ net295 _1656_ _1657_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3459__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2216_ net21 net20 net23 net22 vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3196_ _1391_ _1611_ _1615_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__and3b_1
XFILLER_0_20_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2147_ _0937_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__nor2_4
XFILLER_0_94_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2078_ team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] net110 net134 net764 vssd1
+ vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4719_ net487 vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2976__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output67_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3050_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] _1519_ net200 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[61\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2001_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] net146 net117
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1 vccd1 _0748_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3697__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2805__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3952_ clknet_leaf_34_wb_clk_i _0015_ net268 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2903_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\] net153 _1473_ net785
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[8\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3883_ net283 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2834_ _0515_ _1428_ _1435_ _1411_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2765_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ _1378_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4504_ net315 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3392__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2696_ team_10_WB.instance_to_wrap.message_reg.msg\[4\] team_10_WB.instance_to_wrap.message_reg.msg\[5\]
+ team_10_WB.instance_to_wrap.message_reg.msg\[6\] team_10_WB.instance_to_wrap.message_reg.msg\[7\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4435_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[32\]
+ _0418_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_26_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4366_ clknet_leaf_19_wb_clk_i _0751_ _0349_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3317_ _0815_ net206 _1680_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout290_A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4297_ clknet_leaf_12_wb_clk_i _0687_ _0286_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3248_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\] _1608_ vssd1 vssd1 vccd1
+ vccd1 _1647_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2495__B _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3179_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] _1602_ vssd1 vssd1 vccd1 vccd1
+ _0503_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4565__536 vssd1 vssd1 vccd1 vccd1 net536 _4565__536/LO sky130_fd_sc_hd__conb_1
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2016__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3368__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2949__A2 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2550_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2481_ net598 net132 _1187_ _1213_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4220_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[82\]
+ _0209_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[82\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4151_ clknet_leaf_9_wb_clk_i _0622_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfxtp_2
X_3102_ net200 net684 net187 _1545_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[87\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4082_ clknet_leaf_8_wb_clk_i _0553_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4588__547 vssd1 vssd1 vccd1 vccd1 net547 _4588__547/LO sky130_fd_sc_hd__conb_1
X_3033_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\]
+ net186 vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3935_ net241 vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout136_A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3866_ net282 vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2817_ _0516_ _1409_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3797_ net277 vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2748_ _1369_ _1370_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[17\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout303_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2679_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] _1327_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__a21o_1
X_4671__439 vssd1 vssd1 vccd1 vccd1 _4671__439/HI net439 sky130_fd_sc_hd__conb_1
XFILLER_0_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4418_ clknet_leaf_20_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[15\]
+ _0401_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout301 net303 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4349_ clknet_leaf_14_wb_clk_i _0739_ _0338_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[72\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3356__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2564__B1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1981_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3720_ net234 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ net259 vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2602_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] _1275_ _1285_ net869
+ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3582_ net287 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2533_ net561 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2464_ net734 net128 _1194_ _1205_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4203_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[65\]
+ _0192_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[65\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2395_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked team_10_WB.instance_to_wrap.host_col\[1\]
+ _0850_ _1158_ net648 vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4134_ clknet_leaf_16_wb_clk_i _0605_ _0133_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[69\]
+ sky130_fd_sc_hd__dfrtp_1
X_4065_ clknet_leaf_34_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[2\]
+ _0085_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3016_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\] net184 _1502_ team_10_WB.instance_to_wrap.hostdisp.Cstate
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[44\] sky130_fd_sc_hd__o211a_1
XFILLER_0_91_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout253_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3918_ net242 vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3849_ net254 vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2013__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout120 _1473_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
Xfanout131 _1183_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_4
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_4
Xfanout153 _1182_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4532__343 vssd1 vssd1 vccd1 vccd1 _4532__343/HI net343 sky130_fd_sc_hd__conb_1
Xfanout164 _0872_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2077__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3019__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4693__461 vssd1 vssd1 vccd1 vccd1 _4693__461/HI net461 sky130_fd_sc_hd__conb_1
XANTENNA__2001__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4015__RESET_B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2180_ _0936_ _0961_ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2068__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2473__C1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4752_ net520 vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_2
XFILLER_0_56_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1964_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] net147 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\]
+ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3703_ net233 vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__inv_2
X_4683_ net451 vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1895_ net223 vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3634_ net242 vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3565_ net276 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2516_ net221 _1225_ _1230_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3496_ net276 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__inv_2
X_4516__327 vssd1 vssd1 vccd1 vccd1 _4516__327/HI net327 sky130_fd_sc_hd__conb_1
XFILLER_0_122_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2447_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] net192 vssd1 vssd1 vccd1
+ vccd1 _1197_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2378_ _1130_ _1150_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4117_ clknet_leaf_18_wb_clk_i _0588_ _0116_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4048_ clknet_leaf_7_wb_clk_i _0533_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2059__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4603__377 vssd1 vssd1 vccd1 vccd1 _4603__377/HI net377 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4677__445 vssd1 vssd1 vccd1 vccd1 _4677__445/HI net445 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2959__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1863__A team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4718__486 vssd1 vssd1 vccd1 vccd1 _4718__486/HI net486 sky130_fd_sc_hd__conb_1
XFILLER_0_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold9 team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] vssd1 vssd1 vccd1 vccd1 net561
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2470__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3350_ _1726_ _1729_ net175 vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2301_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] _1078_ _1076_
+ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__o21a_1
XANTENNA__2930__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3281_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ _1664_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2232_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net210 vssd1 vssd1 vccd1
+ vccd1 _1014_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2808__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2163_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2094_ team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] net110 net135 net806 vssd1
+ vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2996_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\] _0838_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ _0839_ net159 vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4735_ net503 vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1947_ net2 _0846_ _0858_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4666_ net434 vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_31_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1878_ net212 vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__inv_2
X_3617_ net246 vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4597_ net197 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3548_ net276 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2921__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3479_ team_10_WB.instance_to_wrap.host_row2\[79\] net165 _1849_ _1851_ vssd1 vssd1
+ vccd1 vccd1 _1852_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2204__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1963__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2912__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3468__A1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2850_ _1444_ _1445_ net174 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2781_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4520_ net331 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_13_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1954__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1954__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4451_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[8\]
+ _0434_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\]
+ sky130_fd_sc_hd__dfstp_1
Xhold206 team_10_WB.instance_to_wrap.dispFSM.guesses\[40\] vssd1 vssd1 vccd1 vccd1
+ net758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\] vssd1 vssd1 vccd1
+ vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold228 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\] vssd1 vssd1 vccd1
+ vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] vssd1 vssd1 vccd1 vccd1
+ net791 sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\] _0815_ net207 _1690_
+ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4382_ clknet_leaf_21_wb_clk_i _0767_ _0365_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2903__B1 _1473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3333_ team_10_WB.instance_to_wrap.host_row1\[40\] _1693_ _1700_ _1712_ vssd1 vssd1
+ vccd1 vccd1 _1713_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3264_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\]
+ _1653_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__and3_2
XFILLER_0_20_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _0997_ _0998_ _0999_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3195_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\] _1390_ vssd1 vssd1 vccd1
+ vccd1 _1615_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2146_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _0939_ _0940_ vssd1 vssd1
+ vccd1 vccd1 _0941_ sky130_fd_sc_hd__or3_2
XFILLER_0_94_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2077_ team_10_WB.instance_to_wrap.dispFSM.guesses\[35\] net111 net136 net870 vssd1
+ vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2979_ _0800_ _1488_ net157 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[21\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3395__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4718_ net486 vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2005__C net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4649_ net417 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2370__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold280_A team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2956__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4609__383 vssd1 vssd1 vccd1 vccd1 _4609__383/HI net383 sky130_fd_sc_hd__conb_1
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3386__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4733__501 vssd1 vssd1 vccd1 vccd1 _4733__501/HI net501 sky130_fd_sc_hd__conb_1
XANTENNA__2212__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4616__387 vssd1 vssd1 vccd1 vccd1 _4616__387/HI net387 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2000_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] net144 net116
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 _0749_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3951_ clknet_leaf_38_wb_clk_i _0014_ net268 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2902_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\] net154 net124 net634
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3882_ net282 vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2833_ _1423_ _1428_ _0518_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3377__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2764_ net843 _1380_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4503_ net314 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_53_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2695_ _1239_ _1246_ _1010_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[2\]
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4434_ clknet_leaf_16_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[31\]
+ _0417_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4365_ clknet_leaf_24_wb_clk_i _0750_ _0348_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[2\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3316_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _1695_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__and3_1
X_4296_ clknet_leaf_15_wb_clk_i _0686_ _0285_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_3247_ _1610_ _1646_ net294 vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3178_ _1277_ _1550_ _1551_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2129_ net133 _0929_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3368__B1 _1746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input11_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2207__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3359__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2480_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] net192 vssd1 vssd1 vccd1
+ vccd1 _1213_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4150_ clknet_leaf_9_wb_clk_i _0621_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
X_3101_ _0788_ net201 vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__nor2_1
X_4081_ clknet_leaf_7_wb_clk_i _0552_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3032_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] _1510_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[52\] sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3934_ net254 vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3865_ net282 vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2816_ _1416_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3796_ net292 vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout129_A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2747_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ _1365_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2678_ net631 _1327_ _1330_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[6\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4417_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[14\]
+ _0400_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4348_ clknet_leaf_31_wb_clk_i net748 _0337_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input3_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4279_ clknet_leaf_29_wb_clk_i _0669_ _0268_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2645__A_N net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1866__A team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1980_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] net144 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3650_ net270 vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2601_ net853 _1275_ _1285_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3581_ net285 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2532_ net610 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2463_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] net195 team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ net125 vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__a22o_1
X_4202_ clknet_leaf_14_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\]
+ _0191_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[64\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2394_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _1089_ _1158_ net659 vssd1
+ vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4133_ clknet_leaf_18_wb_clk_i _0604_ _0132_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ clknet_leaf_35_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[1\]
+ _0084_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3015_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net189 vssd1 vssd1 vccd1
+ vccd1 _1502_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4629__397 vssd1 vssd1 vccd1 vccd1 _4629__397/HI net397 sky130_fd_sc_hd__conb_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout246_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3917_ net250 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3848_ net256 vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3779_ net271 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout110 net111 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__buf_2
Xfanout121 net123 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout132 _1183_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
Xfanout143 _0912_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout165 _1710_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_4
Xfanout176 _1399_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout187 _0994_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
Xfanout198 net63 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1993__C1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2473__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ net519 vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__buf_2
X_1963_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _0874_ _0877_ net158 vssd1
+ vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3702_ net233 vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__inv_2
X_4682_ net450 vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_2
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1894_ team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3633_ net237 vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3564_ net275 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1953__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2515_ net221 _1225_ net191 vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3495_ net236 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__inv_2
X_4555__366 vssd1 vssd1 vccd1 vccd1 _4555__366/HI net366 sky130_fd_sc_hd__conb_1
XFILLER_0_110_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2446_ _1187_ _1196_ net686 net128 vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2377_ _1126_ _1129_ _1128_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout196_A _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4116_ clknet_leaf_17_wb_clk_i _0587_ _0115_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4047_ clknet_leaf_8_wb_clk_i _0532_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3008__A2 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2455__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4498__309 vssd1 vssd1 vccd1 vccd1 _4498__309/HI net309 sky130_fd_sc_hd__conb_1
XFILLER_0_112_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1966__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1981__A2 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2300_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] _1076_ _1077_
+ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3280_ _1666_ _1667_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2231_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] _0803_ vssd1 vssd1 vccd1
+ vccd1 _1013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2162_ _0942_ _0944_ _0956_ net746 vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2093_ team_10_WB.instance_to_wrap.dispFSM.guesses\[19\] net112 net140 net759 vssd1
+ vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2995_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ net159 vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2125__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4734_ net502 vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_2
XFILLER_0_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1946_ _0845_ net194 vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3410__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4665_ net433 vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_114_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1877_ net211 vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3616_ net236 vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__inv_2
X_4596_ net198 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout209_A team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3547_ net277 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4750__518 vssd1 vssd1 vccd1 vccd1 _4750__518/HI net518 sky130_fd_sc_hd__conb_1
XFILLER_0_60_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3478_ team_10_WB.instance_to_wrap.host_row2\[47\] net172 _1708_ team_10_WB.instance_to_wrap.host_row1\[79\]
+ _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2795__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2429_ net628 net130 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\]
+ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__a22o_1
XANTENNA__3477__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2010__D net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__B _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4644__412 vssd1 vssd1 vccd1 vccd1 _4644__412/HI net412 sky130_fd_sc_hd__conb_1
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2988__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1874__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3165__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input41_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3468__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _1390_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4450_ clknet_leaf_25_wb_clk_i net635 _0433_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] vssd1 vssd1 vccd1 vccd1
+ net759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\] vssd1 vssd1 vccd1
+ vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 team_10_WB.instance_to_wrap.dispFSM.guesses\[72\] vssd1 vssd1 vccd1 vccd1
+ net781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3401_ net173 net169 net179 vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__or3_1
X_4381_ clknet_leaf_3_wb_clk_i _0766_ _0364_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_21_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3332_ team_10_WB.instance_to_wrap.host_row1\[72\] _1708_ _1711_ net303 _1706_ vssd1
+ vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_22_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] _1653_ net667 vssd1 vssd1
+ vccd1 vccd1 _1656_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3459__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ net12 net11 net14 net13 vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__or4_4
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3194_ _1390_ _1611_ _1614_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and3b_1
XFILLER_0_20_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2145_ team_10_WB.instance_to_wrap.gamelogic.rights\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2076_ team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] net112 net138 net774 vssd1
+ vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout159_A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2978_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\] net159 _1488_ net210
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[20\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4717_ net485 vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
XANTENNA__3395__B2 team_10_WB.instance_to_wrap.host_row2\[67\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1929_ net223 _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4648_ net416 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4579_ net197 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3083__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3386__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3138__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2212__B net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2897__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 team_10_WB.instance_to_wrap.message_reg.msg\[3\] vssd1 vssd1 vccd1 vccd1 net642
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3950_ clknet_leaf_36_wb_clk_i _0013_ net267 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2901_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\] net151 net122 net708
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[6\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3881_ net282 vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2832_ _1405_ _1433_ _1434_ _1432_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2763_ _1379_ _1380_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[22\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4502_ net313 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2694_ net702 _1009_ _1339_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[1\]
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_129_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4433_ clknet_leaf_17_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[30\]
+ _0416_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_123_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4364_ clknet_leaf_24_wb_clk_i _0749_ _0347_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3315_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ _1682_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2018__C_N net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4295_ clknet_leaf_30_wb_clk_i _0685_ _0284_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_3246_ _1608_ _1645_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3177_ _1283_ _1599_ _1601_ net193 vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2128_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] team_10_WB.instance_to_wrap.buffer.temp_guess\[5\]
+ _0926_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3065__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2059_ net689 net143 net107 net705 vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3368__A1 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4756__524 vssd1 vssd1 vccd1 vccd1 _4756__524/HI net524 sky130_fd_sc_hd__conb_1
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2040__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2207__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4148__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3100_ net205 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] net189 _1544_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[86\] sky130_fd_sc_hd__a31o_1
XFILLER_0_78_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ clknet_leaf_7_wb_clk_i _0551_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3031_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__mux2_1
XANTENNA__2893__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3933_ net270 vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4613__A team_10_WB.instance_to_wrap.blue vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3864_ net287 vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2815_ _0514_ _0515_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3795_ net272 vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2746_ team_10_WB.instance_to_wrap.clock_div.count\[17\] _1367_ vssd1 vssd1 vccd1
+ vccd1 _1369_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2677_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] _1327_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4416_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[13\]
+ _0399_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout303 net6 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_2
X_4571__542 vssd1 vssd1 vccd1 vccd1 net542 _4571__542/LO sky130_fd_sc_hd__conb_1
X_4347_ clknet_leaf_13_wb_clk_i _0737_ _0336_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[70\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4278_ clknet_leaf_30_wb_clk_i _0668_ _0267_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3229_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\]
+ _1632_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\] vssd1 vssd1 vccd1 vccd1
+ _1636_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2261__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1882__A team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2600_ _1270_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3580_ net284 vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2531_ net602 team_10_WB.instance_to_wrap.buffer.temp_guess\[5\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2462_ net564 net129 _1204_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4201_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[63\]
+ _0190_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[63\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2393_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _1093_ _1158_ net655 vssd1
+ vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4132_ clknet_leaf_17_wb_clk_i _0603_ _0131_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4063_ clknet_leaf_35_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[0\]
+ _0083_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3014_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\] net184 _1501_ net205
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\] sky130_fd_sc_hd__o211a_1
XFILLER_0_95_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3916_ net263 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout141_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout239_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3847_ net241 vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3778_ net293 vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2729_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ _1358_ _1177_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout111 _0913_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
Xfanout122 net123 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_4
Xfanout133 _0919_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
Xfanout144 net146 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout155 _1181_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout166 _1710_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
Xfanout177 _1727_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_4
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
Xfanout199 net202 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1877__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2473__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4661__429 vssd1 vssd1 vccd1 vccd1 _4661__429/HI net429 sky130_fd_sc_hd__conb_1
XFILLER_0_5_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4750_ net518 vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__buf_2
XFILLER_0_5_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1962_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] net144 vssd1 vssd1 vccd1
+ vccd1 _0877_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3701_ net231 vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4681_ net449 vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_2
XFILLER_0_28_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1893_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\] vssd1 vssd1 vccd1 vccd1
+ _0817_ sky130_fd_sc_hd__inv_2
XANTENNA__1984__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3632_ net237 vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3563_ net275 vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2514_ _1226_ _1229_ net191 vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__and3b_1
XFILLER_0_122_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3494_ net242 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2445_ _0836_ net192 vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2376_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] _1084_ _1148_
+ _1149_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__o22a_1
X_4115_ clknet_leaf_5_wb_clk_i _0586_ _0114_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout189_A _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ clknet_leaf_7_wb_clk_i _0531_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3413__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3404__B1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2231__A team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2930__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2230_ _0822_ net214 team_10_WB.instance_to_wrap.gamelogic.state\[2\] _0988_ team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__a311o_1
X_2161_ _0942_ _0943_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2092_ team_10_WB.instance_to_wrap.dispFSM.guesses\[20\] net115 net138 net824 vssd1
+ vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2446__B2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2994_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] net157 vssd1 vssd1 vccd1
+ vccd1 _1493_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4733_ net501 vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_2
XFILLER_0_44_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1945_ _0845_ net194 vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__and2_1
X_4522__333 vssd1 vssd1 vccd1 vccd1 _4522__333/HI net333 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1957__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4664_ net432 vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1876_ net210 vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3615_ net237 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4595_ net197 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3546_ net277 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2921__A2 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3477_ team_10_WB.instance_to_wrap.host_row2\[87\] net171 net178 team_10_WB.instance_to_wrap.host_row2\[63\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2428_ net187 _1185_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nand2_1
XANTENNA__2134__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2359_ _1124_ _1134_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4029_ clknet_leaf_6_wb_clk_i _0514_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4683__451 vssd1 vssd1 vccd1 vccd1 _4683__451/HI net451 sky130_fd_sc_hd__conb_1
XFILLER_0_135_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3999__RESET_B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4031__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4724__492 vssd1 vssd1 vccd1 vccd1 _4724__492/HI net492 sky130_fd_sc_hd__conb_1
XFILLER_0_47_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input34_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4506__317 vssd1 vssd1 vccd1 vccd1 _4506__317/HI net317 sky130_fd_sc_hd__conb_1
XFILLER_0_127_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold208 team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] vssd1 vssd1 vccd1 vccd1
+ net760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\] vssd1 vssd1 vccd1
+ vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
X_3400_ _1686_ _1698_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__or3_1
X_4380_ clknet_leaf_23_wb_clk_i _0765_ _0363_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2903__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3331_ team_10_WB.instance_to_wrap.host_row2\[56\] net178 net165 team_10_WB.instance_to_wrap.host_row2\[72\]
+ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ net742 _1653_ _1655_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ net39 net38 net10 net9 vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _1614_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2144_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__a21o_1
X_4667__435 vssd1 vssd1 vccd1 vccd1 _4667__435/HI net435 sky130_fd_sc_hd__conb_1
XFILLER_0_117_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2075_ net673 net141 net107 net685 vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4708__476 vssd1 vssd1 vccd1 vccd1 _4708__476/HI net476 sky130_fd_sc_hd__conb_1
XFILLER_0_18_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2977_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] net162 _1488_ net211
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[19\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1975__A team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3395__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4716_ net484 vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
X_1928_ team_10_WB.instance_to_wrap.host_col\[3\] net222 vssd1 vssd1 vccd1 vccd1 _0851_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_72_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4647_ net415 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4578_ net197 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3529_ net244 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3386__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2594__B1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold80 team_10_WB.instance_to_wrap.host_row1\[40\] vssd1 vssd1 vccd1 vccd1 net632
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] vssd1 vssd1 vccd1
+ vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2900_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\] net154 net124 net574
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3880_ net282 vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2831_ _1430_ _1431_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3377__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2762_ team_10_WB.instance_to_wrap.clock_div.count\[21\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ team_10_WB.instance_to_wrap.clock_div.count\[22\] _1374_ vssd1 vssd1 vccd1 vccd1
+ _1380_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4501_ net312 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2693_ _1009_ _1238_ _1339_ _1340_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[0\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4432_ clknet_leaf_16_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[29\]
+ _0415_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4363_ clknet_leaf_24_wb_clk_i _0748_ _0346_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_26_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3314_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__nand2_2
X_4294_ clknet_leaf_31_wb_clk_i _0684_ _0283_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_3245_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _1645_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3176_ _1582_ _1600_ _0906_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2127_ net133 _0928_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout171_A _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2058_ team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] net114 net138 net797 vssd1
+ vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3359__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XANTENNA_output65_A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_120_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3030_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] _1509_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[51\] sky130_fd_sc_hd__mux2_1
XANTENNA__2893__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3932_ net262 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3863_ net282 vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2814_ _1413_ _1418_ _1416_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3794_ net290 vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2745_ _1367_ _1368_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[16\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2676_ _1318_ _1328_ _1329_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[5\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4415_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[12\]
+ _0398_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4346_ clknet_leaf_28_wb_clk_i net728 _0335_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[69\]
+ sky130_fd_sc_hd__dfrtp_1
X_4277_ clknet_leaf_14_wb_clk_i _0667_ _0266_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3228_ net738 _1633_ _1635_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2089__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3159_ _1586_ _1587_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_42_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2530_ net572 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2461_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] net200 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ _1189_ net128 vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4200_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[62\]
+ _0189_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[62\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2392_ net2 net679 _1158_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4131_ clknet_leaf_10_wb_clk_i _0602_ _0130_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4062_ clknet_leaf_7_wb_clk_i _0547_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3013_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] net190 vssd1 vssd1 vccd1
+ vccd1 _1501_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3915_ net270 vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3440__B2 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3846_ net254 vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3777_ net289 vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2728_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ vssd1 vssd1 vccd1
+ vccd1 _1358_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout301_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2951__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2659_ _1310_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout112 net115 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_4
Xfanout123 _1473_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_2
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4329_ clknet_leaf_12_wb_clk_i _0719_ _0318_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout145 net146 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout156 _0873_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_4
Xfanout167 _1704_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout178 _1709_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_4
Xfanout189 _0994_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2473__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1961_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] net146 net116 net874 vssd1
+ vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__o22a_1
XANTENNA__3422__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3700_ net239 vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__inv_2
X_4680_ net448 vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_2
XFILLER_0_43_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1892_ team_10_WB.instance_to_wrap.lcdPlayer.currentState\[0\] vssd1 vssd1 vccd1
+ vccd1 _0816_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1984__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3631_ net250 vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3562_ net275 vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2933__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2513_ net221 _1225_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] vssd1
+ vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3493_ net236 vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2444_ net597 net132 _1185_ _1195_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2375_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2161__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4114_ clknet_leaf_16_wb_clk_i _0585_ _0113_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4045_ clknet_leaf_7_wb_clk_i _0530_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2139__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2449__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2464__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout251_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3829_ net250 vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1888__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1966__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2915__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2160_ _0936_ _0941_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2091_ team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] net143 net107 net696 vssd1
+ vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2993_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\] net157 _1492_ net208
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[31\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4732_ net500 vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_2
XFILLER_0_127_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1944_ _0858_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4561__372 vssd1 vssd1 vccd1 vccd1 _4561__372/HI net372 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4663_ net431 vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_114_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1875_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1 vccd1
+ _0800_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3614_ net237 vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2422__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4594_ net198 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2906__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3545_ net277 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3108__A_N net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3476_ team_10_WB.instance_to_wrap.host_row1\[55\] _1699_ net167 team_10_WB.instance_to_wrap.host_row1\[63\]
+ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2427_ net183 _1186_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout299_A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3331__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2358_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1133_ _1132_ _1117_
+ _1100_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_100_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2289_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__inv_2
X_4028_ clknet_leaf_10_wb_clk_i _0513_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2437__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input27_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4545__356 vssd1 vssd1 vccd1 vccd1 _4545__356/HI net356 sky130_fd_sc_hd__conb_1
XANTENNA__3389__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2061__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold209 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1 vccd1
+ net761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3010__C1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3330_ _1683_ _1687_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] _1653_ net295 vssd1 vssd1
+ vccd1 vccd1 _1655_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ net19 net8 net33 net30 vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _1389_ _1611_ _1613_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2143_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.correct\[0\]
+ team_10_WB.instance_to_wrap.correct\[2\] vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__o21a_1
X_2074_ team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] net114 net139 net817 vssd1
+ vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2976_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\] net163 _1488_ net212
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[18\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4715_ net483 vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2052__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1927_ net226 _0848_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4646_ net414 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4008__SET_B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4577_ net197 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3528_ net238 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3459_ team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] _1701_ _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3711__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2897__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold70 team_10_WB.instance_to_wrap.host_row1\[56\] vssd1 vssd1 vccd1 vccd1 net622
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] vssd1 vssd1 vccd1
+ vccd1 net633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold92 _0488_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4740__508 vssd1 vssd1 vccd1 vccd1 _4740__508/HI net508 sky130_fd_sc_hd__conb_1
XFILLER_0_15_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2830_ _1430_ _1431_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2761_ net859 _1378_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4500_ net311 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_26_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2692_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] _1241_ vssd1 vssd1
+ vccd1 vccd1 _1340_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4431_ clknet_leaf_17_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[28\]
+ _0414_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4634__402 vssd1 vssd1 vccd1 vccd1 _4634__402/HI net402 sky130_fd_sc_hd__conb_1
XFILLER_0_125_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4362_ clknet_leaf_12_wb_clk_i _0747_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3313_ net206 _1686_ _1688_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__and4b_4
XFILLER_0_21_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4293_ clknet_leaf_13_wb_clk_i _0683_ _0282_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_96_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3244_ _1610_ _1644_ net294 vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3175_ _0887_ _0894_ _0891_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3531__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2126_ net209 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2057_ net722 net142 net108 net745 vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2959_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] _1480_ _1481_ vssd1
+ vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4629_ net397 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3706__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4044__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_78_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3931_ net270 vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3862_ net283 vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2813_ _1415_ _1417_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3793_ net278 vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2744_ team_10_WB.instance_to_wrap.clock_div.count\[16\] _1365_ _1177_ vssd1 vssd1
+ vccd1 vccd1 _1368_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2675_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\]
+ _1321_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\] vssd1 vssd1 vccd1
+ vccd1 _1329_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2430__A _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4414_ clknet_leaf_17_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[11\]
+ _0397_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_26_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4345_ clknet_leaf_13_wb_clk_i _0735_ _0334_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[68\]
+ sky130_fd_sc_hd__dfstp_1
X_4276_ clknet_leaf_48_wb_clk_i _0666_ _0265_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3227_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] _1633_ net170 vssd1
+ vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout281_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3158_ _1560_ _1585_ _1584_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2494__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2109_ team_10_WB.instance_to_wrap.dispFSM.guesses\[3\] net112 net140 net749 vssd1
+ vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__o22a_1
X_3089_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] net195 vssd1 vssd1 vccd1
+ vccd1 _1539_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1996__C1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2460_ net571 net128 _1203_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2391_ net623 _1158_ _1159_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__a21o_1
X_4130_ clknet_leaf_28_wb_clk_i _0601_ _0129_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_4061_ clknet_leaf_7_wb_clk_i _0546_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_3012_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\] net184 _1500_ net203
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[42\] sky130_fd_sc_hd__o211a_1
XFILLER_0_21_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4746__514 vssd1 vssd1 vccd1 vccd1 _4746__514/HI net514 sky130_fd_sc_hd__conb_1
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3914_ net256 vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__inv_2
XANTENNA__2425__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3845_ net247 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3776_ net291 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2727_ _1180_ _1355_ _1357_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[9\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_131_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2951__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2658_ net191 _1234_ _1225_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__o21bai_2
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2589_ _1272_ _1273_ _0902_ _0908_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2703__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_4
Xfanout124 _1472_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_4
X_4328_ clknet_leaf_29_wb_clk_i _0718_ _0317_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[51\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout146 _0862_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input1_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _0873_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
Xfanout168 _1702_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_4
Xfanout179 _1709_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4259_ clknet_leaf_57_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[2\]
+ _0248_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2942__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3407__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1960_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\]
+ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1891_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] vssd1 vssd1 vccd1 vccd1
+ _0815_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3630_ net247 vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3561_ net275 vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2512_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] _1226_ _1228_ vssd1
+ vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3492_ net236 vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2443_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net184 vssd1 vssd1 vccd1
+ vccd1 _1195_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2374_ _0871_ _1147_ _1087_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4113_ clknet_leaf_16_wb_clk_i _0584_ _0112_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4044_ clknet_leaf_7_wb_clk_i _0529_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2449__B1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout244_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3413__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3828_ net262 vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3177__B2 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3759_ net280 vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3714__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2215__D _1000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2090_ team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] net113 net139 net847 vssd1
+ vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2992_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net160 _1491_ team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[30\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ net499 vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1943_ _0844_ _0855_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4662_ net430 vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1874_ net209 vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3613_ net237 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2422__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4593_ net197 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1921__A_N net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3544_ net277 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3475_ team_10_WB.instance_to_wrap.host_row1\[47\] _1693_ _1703_ team_10_WB.instance_to_wrap.host_row1\[71\]
+ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2426_ _0993_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2357_ _0823_ _0828_ _1859_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2288_ team_10_WB.instance_to_wrap.host_col\[3\] net223 team_10_WB.instance_to_wrap.host_col\[0\]
+ net222 vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4027_ clknet_leaf_48_wb_clk_i net567 _0074_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3709__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4651__419 vssd1 vssd1 vccd1 vccd1 _4651__419/HI net419 sky130_fd_sc_hd__conb_1
XFILLER_0_24_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3086__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ net563 _1651_ _1654_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ net35 net34 net37 net36 vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2142_ _0916_ _0935_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2073_ net699 net142 net108 net718 vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3092__A3 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2975_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\] net163 _1488_ net213
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[17\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4714_ net482 vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1926_ net226 _0848_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4645_ net413 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4576_ net198 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3527_ net238 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3458_ team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] net166 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[14\]
+ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2409_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3389_ team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] net171 net179 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\]
+ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3068__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3174__A team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4512__323 vssd1 vssd1 vccd1 vccd1 _4512__323/HI net323 sky130_fd_sc_hd__conb_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold60 team_10_WB.instance_to_wrap.host_row1\[59\] vssd1 vssd1 vccd1 vccd1 net612
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\] vssd1 vssd1 vccd1
+ vccd1 net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[7\] vssd1 vssd1 vccd1 vccd1
+ net634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3059__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold93 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] vssd1 vssd1 vccd1 vccd1
+ net645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4014__SET_B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2760_ _1377_ _1378_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[21\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2691_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] _1246_ _1238_ vssd1
+ vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4430_ clknet_leaf_17_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[27\]
+ _0413_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_2 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4673__441 vssd1 vssd1 vccd1 vccd1 _4673__441/HI net441 sky130_fd_sc_hd__conb_1
X_4361_ clknet_leaf_10_wb_clk_i _0004_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2742__C1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3312_ _1691_ _1692_ net295 vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4292_ clknet_leaf_29_wb_clk_i _0682_ _0281_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3243_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__xnor2_1
X_4714__482 vssd1 vssd1 vccd1 vccd1 _4714__482/HI net482 sky130_fd_sc_hd__conb_1
XFILLER_0_119_1308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3174_ team_10_WB.instance_to_wrap.dispFSM.msg\[6\] _1550_ vssd1 vssd1 vccd1 vccd1
+ _1599_ sky130_fd_sc_hd__or2_1
X_2125_ net133 _0927_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__and2_1
XANTENNA__2428__A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3023__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2056_ team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] net113 net139 net800 vssd1
+ vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2273__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3470__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout157_A _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2958_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] _0832_ net162 vssd1 vssd1 vccd1
+ vccd1 _1481_ sky130_fd_sc_hd__a41o_1
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1909_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\] vssd1 vssd1 vccd1 vccd1
+ _0832_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2889_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] net1 _1469_ vssd1 vssd1 vccd1
+ vccd1 _1470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4628_ net396 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XFILLER_0_128_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4559_ net370 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3722__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3461__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4657__425 vssd1 vssd1 vccd1 vccd1 _4657__425/HI net425 sky130_fd_sc_hd__conb_1
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2801__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_120_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_78_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3930_ net257 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3452__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3861_ net283 vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2812_ _0816_ _0817_ net176 vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3792_ net289 vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2743_ team_10_WB.instance_to_wrap.clock_div.count\[15\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ _1364_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2674_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4413_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[10\]
+ _0396_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_125_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2430__B _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4344_ clknet_leaf_28_wb_clk_i _0734_ _0333_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[67\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4275_ clknet_leaf_48_wb_clk_i _0665_ _0264_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3226_ net865 _1632_ _1634_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3157_ _1560_ _1584_ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout274_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2108_ team_10_WB.instance_to_wrap.dispFSM.guesses\[4\] net114 net138 net840 vssd1
+ vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__o22a_1
X_3088_ net199 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] net185 _1538_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[80\] sky130_fd_sc_hd__a31o_1
XFILLER_0_136_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2039_ team_10_WB.instance_to_wrap.dispFSM.guesses\[73\] net109 net135 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__o22a_1
XANTENNA__3443__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2246__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3717__A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2237__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2390_ _0858_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__nor2_1
XANTENNA_output70_A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4060_ clknet_leaf_7_wb_clk_i _0545_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3011_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] net190 vssd1 vssd1 vccd1
+ vccd1 _1500_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3425__B1 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3913_ net258 vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2425__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1987__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3844_ net262 vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3775_ net280 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__inv_2
XANTENNA__3537__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2726_ _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2657_ net191 _1225_ _1227_ _1234_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[2\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2588_ _0898_ _0901_ _0907_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4327_ clknet_leaf_29_wb_clk_i _0717_ _0316_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[50\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout114 net115 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_4
Xfanout125 _1191_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_4
XANTENNA__3272__A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout136 _0914_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout158 _0873_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_4
X_4258_ clknet_leaf_56_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[1\]
+ _0247_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout169 _1702_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3209_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] _1621_ _1623_ vssd1 vssd1
+ vccd1 vccd1 _0535_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4189_ clknet_leaf_19_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[51\]
+ _0178_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[51\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3416__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1978__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1890_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ _0814_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3560_ net275 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__inv_2
XANTENNA__2933__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2511_ _1225_ _1227_ net191 vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3491_ net242 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2442_ net609 net129 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\]
+ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3343__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2373_ _1137_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4112_ clknet_leaf_27_wb_clk_i net617 _0111_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4043_ clknet_leaf_7_wb_clk_i _0528_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3031__S net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3827_ net247 vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3758_ net291 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2709_ _1345_ _1346_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
X_3689_ net231 vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2612__A1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2915__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2128__A0 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2991_ net710 net157 _1492_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[29\] sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4730_ net498 vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1942_ _0819_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4661_ net429 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_127_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1873_ net208 vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3612_ net285 vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4592_ net551 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2906__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3543_ net279 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3474_ team_10_WB.instance_to_wrap.dispFSM.guesses\[31\] net169 net166 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\]
+ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2425_ net196 _0942_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3026__S net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3331__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2356_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1119_ vssd1 vssd1 vccd1
+ vccd1 _1132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2287_ _1064_ _1063_ team_10_WB.instance_to_wrap.gamelogic.rights\[0\] vssd1 vssd1
+ vccd1 vccd1 _0644_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout187_A _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4026_ clknet_leaf_48_wb_clk_i net573 _0073_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4568__539 vssd1 vssd1 vccd1 vccd1 net539 _4568__539/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4690__458 vssd1 vssd1 vccd1 vccd1 _4690__458/HI net458 sky130_fd_sc_hd__conb_1
XFILLER_0_63_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4731__499 vssd1 vssd1 vccd1 vccd1 _4731__499/HI net499 sky130_fd_sc_hd__conb_1
XFILLER_0_76_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3389__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2061__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _0806_ _0996_ net192 _0945_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ net576 _1612_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2141_ _0916_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2072_ team_10_WB.instance_to_wrap.dispFSM.guesses\[40\] net112 net140 net825 vssd1
+ vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2974_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] net163 _1488_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[16\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_4713_ net481 vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
X_1925_ net2 net3 net300 vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_45_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4644_ net412 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4575_ net198 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3526_ net238 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3457_ team_10_WB.instance_to_wrap.host_row1\[78\] _1708_ _1829_ _1830_ vssd1 vssd1
+ vccd1 vccd1 _1831_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2408_ _1164_ _1167_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__nor3_1
X_3388_ team_10_WB.instance_to_wrap.dispFSM.guesses\[75\] _1715_ _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[11\]
+ _1764_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__a221o_1
X_2339_ _1110_ _1111_ _1113_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4009_ clknet_leaf_32_wb_clk_i _0497_ net271 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input32_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4551__362 vssd1 vssd1 vccd1 vccd1 _4551__362/HI net362 sky130_fd_sc_hd__conb_1
Xhold50 team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] vssd1 vssd1 vccd1 vccd1 net602
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 team_10_WB.instance_to_wrap.host_row1\[57\] vssd1 vssd1 vccd1 vccd1 net613
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] vssd1 vssd1 vccd1
+ vccd1 net624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[7\] vssd1 vssd1 vccd1
+ vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2253__B net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2690_ net784 _1336_ _1338_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_3 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4360_ clknet_leaf_10_wb_clk_i _0003_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3311_ net176 net683 vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__nand2b_1
X_4291_ clknet_leaf_13_wb_clk_i _0681_ _0280_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3242_ net646 _1610_ net293 vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__a21oi_1
X_3173_ _0903_ _1298_ _1598_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2124_ net208 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0927_ sky130_fd_sc_hd__mux2_1
XANTENNA__2428__B _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2055_ team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] net109 net135 team_10_WB.instance_to_wrap.dispFSM.guesses\[65\]
+ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2273__A2 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2957_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] _0833_ net161 vssd1 vssd1 vccd1
+ vccd1 _1480_ sky130_fd_sc_hd__a41o_1
XFILLER_0_106_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1908_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1 vssd1 vccd1 vccd1
+ _0831_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2888_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] vssd1 vssd1 vccd1 vccd1
+ _1469_ sky130_fd_sc_hd__and3b_1
XANTENNA__2981__A0 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4627_ net395 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_114_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4494__305 vssd1 vssd1 vccd1 vccd1 _4494__305/HI net305 sky130_fd_sc_hd__conb_1
XFILLER_0_13_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4558_ net369 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_114_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3509_ net236 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__inv_2
X_4489_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[46\]
+ _0472_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4535__346 vssd1 vssd1 vccd1 vccd1 _4535__346/HI net346 sky130_fd_sc_hd__conb_1
XFILLER_0_25_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4696__464 vssd1 vssd1 vccd1 vccd1 _4696__464/HI net464 sky130_fd_sc_hd__conb_1
XFILLER_0_23_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_128_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_0_37_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4090__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3860_ net287 vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2811_ _1413_ _1415_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3791_ net280 vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2742_ net829 _1364_ _1366_ _1177_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[15\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2673_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ _1324_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4412_ clknet_leaf_16_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[9\]
+ _0395_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4343_ clknet_leaf_29_wb_clk_i _0733_ _0332_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[66\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4274_ clknet_leaf_48_wb_clk_i _0664_ _0263_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3225_ net170 _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3156_ _1569_ _1574_ _1573_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2107_ net698 net141 net107 net709 vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3087_ _0790_ net199 vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2038_ team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] net111 net136 net838 vssd1
+ vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__o22a_1
XFILLER_0_136_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3989_ clknet_leaf_53_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[26\]
+ _0057_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2954__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1996__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3908__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3370__B1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_output63_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3010_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\] net183 _1499_ net199
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[41\] sky130_fd_sc_hd__o211a_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3912_ net257 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3843_ net247 vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3774_ net289 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2936__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2725_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ team_10_WB.instance_to_wrap.clock_div.count\[9\] _1351_ vssd1 vssd1 vccd1 vccd1
+ _1356_ sky130_fd_sc_hd__and4_2
XANTENNA__3029__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2656_ _1307_ _1316_ _1314_ _1228_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[1\]
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2587_ net5 _0902_ _0904_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_41_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2164__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3361__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4326_ clknet_leaf_30_wb_clk_i _0716_ _0315_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[49\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout115 _0913_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_2
Xfanout126 _1188_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
Xfanout137 net139 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xfanout148 _0862_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_4
Xfanout159 net164 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_4257_ clknet_leaf_57_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[0\]
+ _0246_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3208_ net170 _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__nor2_1
X_4188_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[50\]
+ _0177_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[50\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2467__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3139_ _1286_ _1554_ _1565_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2927__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold180 _1387_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3352__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] vssd1 vssd1 vccd1 vccd1
+ net743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3407__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1969__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1969__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2510_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net221 vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3490_ net247 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4752__520 vssd1 vssd1 vccd1 vccd1 _4752__520/HI net520 sky130_fd_sc_hd__conb_1
XFILLER_0_110_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2441_ net669 net130 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\]
+ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3343__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2372_ _1131_ _1135_ _1096_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4111_ clknet_leaf_10_wb_clk_i net707 _0110_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4042_ clknet_leaf_7_wb_clk_i _0527_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout132_A _1183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3826_ net258 vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2909__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3757_ net278 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2385__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2708_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ net836 vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3688_ net231 vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2639_ _0946_ _1304_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[0\]
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4309_ clknet_leaf_14_wb_clk_i _0699_ _0298_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_76_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4151__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4736__504 vssd1 vssd1 vccd1 vccd1 _4736__504/HI net504 sky130_fd_sc_hd__conb_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3325__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3921__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2256__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2990_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] net161 _1491_ net210
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[28\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1941_ net226 _0848_ _0851_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4660_ net428 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1872_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1 vccd1
+ _0797_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3087__B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3611_ net249 vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4591_ net550 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XANTENNA__2367__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3542_ net239 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3473_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] net167 _1844_ _1845_ vssd1 vssd1
+ vccd1 vccd1 _1846_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2424_ net196 _0942_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__nor2_4
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2355_ _1128_ _1129_ _1126_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_23_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2286_ _0940_ _1064_ _1065_ _1063_ net798 vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4025_ clknet_leaf_48_wb_clk_i net603 _0072_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3042__S net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3809_ net273 vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3010__A2 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2140_ _0822_ team_10_WB.instance_to_wrap.gamelogic.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2071_ team_10_WB.instance_to_wrap.dispFSM.guesses\[41\] net110 net134 net835 vssd1
+ vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2037__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2973_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] net125 _1486_ _1487_
+ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__nand4_4
XFILLER_0_45_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4712_ net480 vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
XFILLER_0_127_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1924_ net299 net3 vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4643_ net411 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_115_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4574_ net198 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3525_ net230 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3037__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3456_ team_10_WB.instance_to_wrap.host_row1\[46\] _1693_ net172 team_10_WB.instance_to_wrap.host_row2\[46\]
+ _1826_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2407_ _1168_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__or2_1
X_3387_ team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] net166 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2338_ _0811_ _1093_ _1107_ _1108_ _1109_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2269_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net209 vssd1 vssd1 vccd1
+ vccd1 _1051_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4008_ clknet_leaf_32_wb_clk_i _0496_ net273 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold40 team_10_WB.instance_to_wrap.host_row1\[53\] vssd1 vssd1 vccd1 vccd1 net592
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _0510_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_10_WB.instance_to_wrap.host_row1\[52\] vssd1 vssd1 vccd1 vccd1 net614
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_10_WB.instance_to_wrap.host_row1\[41\] vssd1 vssd1 vccd1 vccd1 net636
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] vssd1 vssd1 vccd1
+ vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_45_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2990__B2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 _1003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3310_ _1684_ _1689_ _1690_ net175 vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__or4b_1
XFILLER_0_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4290_ clknet_leaf_29_wb_clk_i _0680_ _0279_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3241_ net587 _1642_ _1643_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3172_ _1290_ _1597_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] vssd1 vssd1 vccd1
+ vccd1 _1598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2123_ _0918_ _0925_ _0922_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2054_ team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] net109 net134 net778 vssd1
+ vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3470__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4641__409 vssd1 vssd1 vccd1 vccd1 _4641__409/HI net409 sky130_fd_sc_hd__conb_1
XFILLER_0_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2956_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\] net156 vssd1 vssd1 vccd1
+ vccd1 _1479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1907_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] vssd1 vssd1 vccd1 vccd1
+ _0830_ sky130_fd_sc_hd__inv_2
X_2887_ net191 _1468_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[5\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_114_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3556__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4626_ net394 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_60_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4557_ net368 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3508_ net235 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4488_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[45\]
+ _0471_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3439_ team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.dispFSM.guesses\[5\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__mux2_1
XANTENNA__3291__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2497__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2249__B1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3461__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_102_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput63 net198 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_101_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3452__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2810_ _1415_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3790_ net291 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2741_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2963__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2672_ net627 _1324_ _1326_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3095__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4411_ clknet_leaf_16_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[8\]
+ _0394_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_125_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4558__369 vssd1 vssd1 vccd1 vccd1 _4558__369/HI net369 sky130_fd_sc_hd__conb_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4342_ clknet_leaf_31_wb_clk_i _0732_ _0331_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[65\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4273_ clknet_leaf_49_wb_clk_i _0663_ _0262_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3224_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1632_ vssd1 vssd1 vccd1
+ vccd1 _1633_ sky130_fd_sc_hd__and2_1
.ends

