* NGSPICE file created from team_11_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt team_11_Wrapper gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36] gpio_in[37] gpio_in[3] gpio_in[4]
+ gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10]
+ gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17]
+ gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23]
+ gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2]
+ gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34] gpio_oeb[35] gpio_oeb[36]
+ gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8]
+ gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14]
+ gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20]
+ gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27]
+ gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33]
+ gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3] gpio_out[4] gpio_out[5]
+ gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1] irq[2] vccd1 vssd1
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__1725__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1270_ net275 _0230_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0985_ net376 net103 net82 _0611_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1606_ clknet_leaf_18_wb_clk_i _0120_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[106\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout127 net134 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_2
Xfanout105 net108 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_4
Xfanout116 _0588_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dlymetal6s2s_1
X_1537_ clknet_leaf_8_wb_clk_i _0051_ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[37\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_2
X_1468_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[37\] _0342_ _0347_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[29\] vssd1 vssd1 vccd1
+ vccd1 _0407_ sky130_fd_sc_hd__a22o_1
X_1399_ net118 net93 _0318_ _0320_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__and4_4
XTAP_TAPCELL_ROW_38_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1427__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold122_A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ _0465_ _0466_ _0470_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1322_ _0020_ _0581_ net187 _0479_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__and4b_1
X_1253_ net294 _0539_ _0222_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__o21a_1
X_1184_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[117\] net143 net125
+ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0968_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\] net145 net122
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[25\] net95 vssd1 vssd1
+ vccd1 vccd1 _0603_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout125_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0899_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[5\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[4\]
+ _0547_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1345__A0 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1441__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0822_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[11\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[10\]
+ _0498_ _0501_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0753_ net270 net39 _0456_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1305_ _0582_ _0237_ _0260_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__o21ai_2
X_1236_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[4\] net307 net186 vssd1
+ vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1167_ net336 net103 net82 _0702_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1098_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[74\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[90\] net99 vssd1 vssd1
+ vccd1 vccd1 _0668_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1021_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[43\] net112 _0629_
+ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__o21a_1
X_1760__255 vssd1 vssd1 vccd1 vccd1 net255 _1760__255/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_45_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1785_ net208 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_21_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0805_ net323 _0494_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0736_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[29\] vssd1 vssd1 vccd1 vccd1
+ _0442_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1219_ team_11_WB.instance_to_wrap.sending.currentState\[0\] team_11_WB.instance_to_wrap.sending.currentState\[1\]
+ team_11_WB.instance_to_wrap.sending.currentState\[2\] team_11_WB.instance_to_wrap.sending.currentState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_23_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold30 team_11_WB.instance_to_wrap.sending.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[13\] vssd1 vssd1 vccd1 vccd1
+ net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[17\] vssd1 vssd1 vccd1 vccd1
+ net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[21\] vssd1 vssd1 vccd1 vccd1
+ net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[4\] vssd1 vssd1 vccd1 vccd1
+ net323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold96 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[20\] vssd1 vssd1
+ vccd1 vccd1 net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[90\] vssd1 vssd1
+ vccd1 vccd1 net345 sky130_fd_sc_hd__dlygate4sd3_1
X_1744__239 vssd1 vssd1 vccd1 vccd1 net239 _1744__239/LO sky130_fd_sc_hd__conb_1
XFILLER_0_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1490__A2 _0342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1570_ clknet_leaf_13_wb_clk_i _0084_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1004_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[27\] net147 net130
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[43\] net98 vssd1 vssd1
+ vccd1 vccd1 _0621_ sky130_fd_sc_hd__a221o_1
XANTENNA__1481__A2 _0336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1837_ net155 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1768_ net195 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1699_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[14\]
+ net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1472__A2 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__clkbuf_4
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1463__A2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1622_ clknet_leaf_19_wb_clk_i _0136_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1553_ clknet_leaf_8_wb_clk_i _0067_ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[53\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1484_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[38\] _0342_ _0347_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[30\] _0417_ vssd1 vssd1
+ vccd1 vccd1 _0422_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1815__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1445__A2 _0342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0956__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1436__A2 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0984_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[17\] net144 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[33\] vssd1 vssd1 vccd1
+ vccd1 _0611_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1605_ clknet_leaf_21_wb_clk_i _0119_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_1536_ clknet_leaf_26_wb_clk_i _0050_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[36\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout117 _0541_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_2
Xfanout128 net134 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_2
Xfanout106 net108 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_2
Xfanout139 net151 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dlymetal6s2s_1
X_1467_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[45\] _0336_ _0344_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[85\] vssd1 vssd1 vccd1
+ vccd1 _0406_ sky130_fd_sc_hd__a22o_1
X_1398_ net118 net93 _0215_ _0322_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__and4_4
XTAP_TAPCELL_ROW_38_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1427__A2 _0346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1363__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1687__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1321_ net187 _0248_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nand2_1
X_1252_ _0540_ _0535_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__nand2b_1
X_1183_ net319 net103 net82 _0710_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1409__A2 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0967_ net340 net107 _0602_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0898_ _0541_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1519_ clknet_leaf_17_wb_clk_i _0033_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1033__B1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0821_ net337 _0502_ _0505_ _0491_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[10\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0752_ net40 net38 net41 _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1304_ net152 _0587_ _0254_ _0259_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__or4_2
XFILLER_0_36_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1235_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[3\] net303 net186 vssd1
+ vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1166_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[108\] net137 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[124\] vssd1 vssd1 vccd1
+ vccd1 _0702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1097_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[81\] net109 net85
+ _0667_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1015__B1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1823__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1631__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1020_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[35\] net147 net130
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[51\] net99 vssd1 vssd1
+ vccd1 vccd1 _0629_ sky130_fd_sc_hd__a221o_1
XANTENNA__1493__B1 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0804_ _0494_ _0495_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
X_1784_ net207 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_52_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0735_ net187 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout185_A team_11_WB.instance_to_wrap.kp.buffertop.nrst vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1218_ team_11_WB.instance_to_wrap.sending.currentState\[0\] team_11_WB.instance_to_wrap.sending.currentState\[1\]
+ team_11_WB.instance_to_wrap.sending.currentState\[2\] vssd1 vssd1 vccd1 vccd1 _0205_
+ sky130_fd_sc_hd__nor3b_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1149_ net367 net115 net88 _0693_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__o22a_1
XANTENNA__1484__B1 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout98_A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[24\] vssd1 vssd1 vccd1 vccd1
+ net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[23\] vssd1 vssd1 vccd1 vccd1
+ net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[12\] vssd1 vssd1 vccd1 vccd1
+ net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 net42 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[121\] vssd1 vssd1
+ vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[82\] vssd1 vssd1
+ vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[74\] vssd1 vssd1
+ vccd1 vccd1 net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[110\] vssd1 vssd1
+ vccd1 vccd1 net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1003_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[34\] net111 net86
+ _0620_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1466__B1 _0349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1836_ net155 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1767_ net194 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1698_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[13\]
+ net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1457__B1 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
Xoutput76 net153 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1448__B1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1621_ clknet_leaf_21_wb_clk_i _0135_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1552_ clknet_leaf_26_wb_clk_i _0066_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1483_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[110\] _0338_ _0340_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[6\] _0420_ vssd1 vssd1
+ vccd1 vccd1 _0421_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1439__B1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout148_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1773__200 vssd1 vssd1 vccd1 vccd1 _1773__200/HI net200 sky130_fd_sc_hd__conb_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1819_ net155 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780__259 vssd1 vssd1 vccd1 vccd1 net259 _1780__259/LO sky130_fd_sc_hd__conb_1
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1217__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0983_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[24\] net107 _0610_
+ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1604_ clknet_leaf_24_wb_clk_i _0118_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1535_ clknet_leaf_18_wb_clk_i _0049_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[35\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout129 net134 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
Xfanout107 net108 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_2
Xfanout118 _0724_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_2
X_1466_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[101\] _0343_ _0349_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[21\] vssd1 vssd1 vccd1
+ vccd1 _0405_ sky130_fd_sc_hd__a22o_1
X_1397_ _0210_ _0317_ _0318_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__and3_4
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1826__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1320_ net187 _0479_ _0581_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__and3_1
X_1251_ _0539_ _0221_ net117 vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__o21bai_1
X_1182_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[116\] net137 vssd1
+ vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_20_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0966_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[8\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[24\] net97 vssd1 vssd1
+ vccd1 vccd1 _0602_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_9_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0897_ _0548_ _0552_ _0553_ _0554_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__or4_4
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1518_ clknet_leaf_19_wb_clk_i _0032_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1449_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[99\] _0343_ _0350_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[59\] vssd1 vssd1 vccd1
+ vccd1 _0390_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0820_ _0504_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0751_ net153 vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1303_ net152 _0587_ _0254_ _0259_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__nor4_2
X_1234_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[2\] net306 net186 vssd1
+ vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__mux2_1
X_1165_ net326 net115 net88 _0701_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_48_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1096_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[73\] net144 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[89\] vssd1 vssd1 vccd1
+ vccd1 _0667_ sky130_fd_sc_hd__a22o_1
XANTENNA__1507__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout130_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0949_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[0\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[16\] vssd1 vssd1 vccd1
+ vccd1 _0593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0803_ net282 _0492_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__nor2_1
X_1783_ net206 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0734_ team_11_WB.instance_to_wrap.sending.currentState\[5\] vssd1 vssd1 vccd1 vccd1
+ _0440_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1181__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1217_ team_11_WB.instance_to_wrap.sending.currentState\[2\] _0204_ net135 vssd1
+ vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout178_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1148_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[99\] net150 net133
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[115\] vssd1 vssd1 vccd1
+ vccd1 _0693_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1079_ net395 net105 net83 _0658_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold21 team_11_WB.instance_to_wrap.sending.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1
+ net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 team_11_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[5\] vssd1 vssd1
+ vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_11_WB.instance_to_wrap.sending.cnt_500hz\[7\] vssd1 vssd1 vccd1 vccd1
+ net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[3\] vssd1 vssd1
+ vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[2\] vssd1 vssd1 vccd1 vccd1
+ net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[49\] vssd1 vssd1
+ vccd1 vccd1 net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[60\] vssd1 vssd1
+ vccd1 vccd1 net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[116\] vssd1 vssd1
+ vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_1002_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[26\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[42\] vssd1 vssd1 vccd1
+ vccd1 _0620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1835_ net154 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1766_ net193 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1697_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[12\]
+ net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1750__245 vssd1 vssd1 vccd1 vccd1 net245 _1750__245/LO sky130_fd_sc_hd__conb_1
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XANTENNA_input23_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1448__B2 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1620_ clknet_leaf_2_wb_clk_i _0134_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1551_ clknet_leaf_18_wb_clk_i _0065_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_1482_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[54\] _0339_ _0341_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[126\] vssd1 vssd1 vccd1
+ vccd1 _0420_ sky130_fd_sc_hd__a22o_1
XANTENNA__1136__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1818_ net232 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1814__231 vssd1 vssd1 vccd1 vccd1 _1814__231/HI net231 sky130_fd_sc_hd__conb_1
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1749_ net244 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1703__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0982_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[16\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[32\] net97 vssd1 vssd1
+ vccd1 vccd1 _0610_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1603_ clknet_leaf_23_wb_clk_i _0117_ net169 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1534_ clknet_leaf_21_wb_clk_i _0048_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout119 net126 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_2
Xfanout108 _0588_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
X_1465_ net267 net135 net167 _0404_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__o211a_1
X_1396_ _0210_ _0215_ _0317_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_38_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout160_A team_11_WB.instance_to_wrap.kp.buffertop.nrst vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold140 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[108\] vssd1 vssd1
+ vccd1 vccd1 net400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1696__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1756__251 vssd1 vssd1 vccd1 vccd1 net251 _1756__251/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_58_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1228__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1250_ net338 _0538_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__nor2_1
X_1181_ net311 net115 net88 _0709_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0965_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[15\] net102 _0601_
+ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0896_ _0548_ _0552_ _0553_ _0554_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__nor4_4
XFILLER_0_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1517_ clknet_leaf_23_wb_clk_i _0031_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1448_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[51\] _0339_ _0340_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[3\] vssd1 vssd1 vccd1 vccd1
+ _0389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1379_ net272 _0557_ _0327_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_2_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1018__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1837__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout90 _0263_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
XFILLER_0_37_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0750_ _0449_ _0450_ _0451_ _0454_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__or4_1
XFILLER_0_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1302_ _0238_ _0241_ _0244_ _0258_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__or4_2
X_1233_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[1\] net304 net186 vssd1
+ vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__mux2_1
X_1164_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[107\] net150 net133
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[123\] vssd1 vssd1 vccd1
+ vccd1 _0701_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1095_ net397 net105 net83 _0666_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0948_ net96 _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0879_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[1\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1493__A2 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0802_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[1\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[0\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[3\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__and4_1
X_1782_ net205 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0733_ team_11_WB.instance_to_wrap.sending.currentState\[2\] vssd1 vssd1 vccd1 vccd1
+ _0439_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1216_ _0202_ _0203_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__and2_1
X_1147_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[106\] net111 net86
+ _0692_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__o22a_1
XANTENNA__1728__RESET_B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1484__A2 _0342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1078_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[64\] net142 net124
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[80\] vssd1 vssd1 vccd1
+ vccd1 _0658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold11 team_11_WB.instance_to_wrap.sending.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[3\] vssd1 vssd1 vccd1 vccd1
+ net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[6\] vssd1 vssd1
+ vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[1\] vssd1 vssd1
+ vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[1\] vssd1 vssd1 vccd1 vccd1
+ net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[10\] vssd1 vssd1 vccd1 vccd1
+ net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[36\] vssd1 vssd1
+ vccd1 vccd1 net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[115\] vssd1 vssd1
+ vccd1 vccd1 net326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[88\] vssd1 vssd1
+ vccd1 vccd1 net359 sky130_fd_sc_hd__dlygate4sd3_1
X_1824__233 vssd1 vssd1 vccd1 vccd1 _1824__233/HI net233 sky130_fd_sc_hd__conb_1
XANTENNA__1475__A2 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1764__191 vssd1 vssd1 vccd1 vccd1 _1764__191/HI net191 sky130_fd_sc_hd__conb_1
X_1001_ net363 net103 _0619_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1466__A2 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1834_ net237 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1765_ net192 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1696_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[11\]
+ net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1808__228 vssd1 vssd1 vccd1 vccd1 _1808__228/HI net228 sky130_fd_sc_hd__conb_1
XANTENNA__1457__A2 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0968__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1448__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0959__A1 team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1550_ clknet_leaf_20_wb_clk_i _0064_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1481_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[46\] _0336_ _0345_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[70\] _0418_ vssd1 vssd1
+ vccd1 vccd1 _0419_ sky130_fd_sc_hd__a221o_1
XANTENNA__1439__A2 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1817_ net154 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1748_ net243 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
X_1679_ clknet_leaf_0_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[3\]
+ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input8_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0981_ net380 net102 _0609_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1602_ clknet_leaf_13_wb_clk_i _0116_ net183 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1533_ clknet_leaf_23_wb_clk_i _0047_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1464_ _0399_ _0400_ _0401_ _0403_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__or4_1
Xfanout109 net116 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1395_ _0199_ _0215_ _0335_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__and3_4
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout153_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold130 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[111\] vssd1 vssd1
+ vccd1 vccd1 net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[46\] vssd1 vssd1
+ vccd1 vccd1 net401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[115\] net150 vssd1
+ vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0964_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[7\] net139 net120
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[23\] net96 vssd1 vssd1
+ vccd1 vccd1 _0601_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0895_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[13\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _0555_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1516_ clknet_leaf_16_wb_clk_i _0030_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1447_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[67\] _0345_ _0349_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[19\] _0387_ vssd1 vssd1
+ vccd1 vccd1 _0388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1378_ net94 _0212_ _0320_ _0323_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__a311o_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1793__216 vssd1 vssd1 vccd1 vccd1 _1793__216/HI net216 sky130_fd_sc_hd__conb_1
XFILLER_0_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout91 _0598_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_2
XFILLER_0_36_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1301_ _0216_ _0237_ _0240_ _0584_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__a31oi_1
X_1232_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[0\] net286 net186 vssd1
+ vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__mux2_1
X_1163_ net387 net111 net86 _0700_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1094_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[72\] net140 net124
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[88\] vssd1 vssd1 vccd1
+ vccd1 _0666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0947_ _0459_ _0590_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0878_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[1\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0752__A net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1411__B1 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1801__223 vssd1 vssd1 vccd1 vccd1 _1801__223/HI net223 sky130_fd_sc_hd__conb_1
X_1781_ net260 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_0_21_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1477__B _0556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0801_ _0492_ _0493_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0732_ team_11_WB.instance_to_wrap.sending.currentState\[1\] vssd1 vssd1 vccd1 vccd1
+ _0438_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1469__B1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1215_ team_11_WB.instance_to_wrap.sending.currentState\[5\] _0716_ _0201_ team_11_WB.instance_to_wrap.sending.currentState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1146_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[98\] net147 net130
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[114\] vssd1 vssd1 vccd1
+ vccd1 _0692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1077_ net377 net110 _0657_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold12 team_11_WB.instance_to_wrap.sending.lcd_rs vssd1 vssd1 vccd1 vccd1 net272
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[7\] vssd1 vssd1
+ vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 team_11_WB.instance_to_wrap.sending.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[122\] vssd1 vssd1
+ vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[1\] vssd1 vssd1 vccd1
+ vccd1 net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_11_WB.instance_to_wrap.sending.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1
+ net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 team_11_WB.instance_to_wrap.sending.cnt_20ms\[4\] vssd1 vssd1 vccd1 vccd1
+ net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[56\] vssd1 vssd1
+ vccd1 vccd1 net349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1000_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[25\] net137 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[41\] net95 vssd1 vssd1
+ vccd1 vccd1 _0619_ sky130_fd_sc_hd__a221o_1
X_1799__222 vssd1 vssd1 vccd1 vccd1 _1799__222/HI net222 sky130_fd_sc_hd__conb_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1833_ net154 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1764_ net191 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1695_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[10\]
+ net161 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout183_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1129_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[97\] net109 _0683_
+ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1531__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XANTENNA_fanout96_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_59_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_1_1__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1619__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1480_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[86\] _0344_ _0351_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[94\] vssd1 vssd1 vccd1
+ vccd1 _0418_ sky130_fd_sc_hd__a22o_1
XANTENNA__1136__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1816_ net154 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1747_ net242 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_1678_ clknet_leaf_0_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[2\]
+ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1712__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[15\] net136 net120
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[31\] net96 vssd1 vssd1
+ vccd1 vccd1 _0609_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1601_ clknet_leaf_10_wb_clk_i _0115_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[101\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_35_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1532_ clknet_leaf_16_wb_clk_i _0046_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1463_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[124\] _0341_ _0344_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[84\] _0402_ vssd1 vssd1
+ vccd1 vccd1 _0403_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1394_ net93 _0318_ _0321_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__and3_4
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout146_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold120 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[23\] vssd1 vssd1
+ vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[91\] vssd1 vssd1
+ vccd1 vccd1 net402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[99\] vssd1 vssd1
+ vccd1 vccd1 net391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0963_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\] net115 net88
+ _0600_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__o22a_1
X_0894_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[5\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[7\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[6\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__or4b_2
XFILLER_0_55_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1515_ clknet_leaf_24_wb_clk_i _0029_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1446_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[123\] _0341_ _0348_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[75\] vssd1 vssd1 vccd1
+ vccd1 _0387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1377_ _0199_ _0212_ _0321_ _0325_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout92 _0598_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1300_ _0584_ _0237_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__nor2_1
X_1231_ team_11_WB.instance_to_wrap.sending.currentState\[5\] _0215_ _0556_ vssd1
+ vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__mux2_1
X_1162_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[106\] net147 net130
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[122\] vssd1 vssd1 vccd1
+ vccd1 _0700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ net362 net110 _0665_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0946_ _0001_ _0020_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__or2_2
X_0877_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[0\] net117 vssd1 vssd1 vccd1
+ vccd1 _0003_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1429_ _0367_ _0368_ _0369_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__or4_1
X_1746__241 vssd1 vssd1 vccd1 vccd1 net241 _1746__241/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_26_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input39_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0943__A team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0800_ net409 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[0\] net314 vssd1 vssd1
+ vccd1 vccd1 _0493_ sky130_fd_sc_hd__a21oi_1
X_1780_ net259 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
X_0731_ team_11_WB.instance_to_wrap.sending.currentState\[0\] vssd1 vssd1 vccd1 vccd1
+ _0437_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1214_ team_11_WB.instance_to_wrap.sending.currentState\[4\] team_11_WB.instance_to_wrap.sending.currentState\[5\]
+ _0717_ team_11_WB.instance_to_wrap.sending.currentState\[0\] _0438_ vssd1 vssd1
+ vccd1 vccd1 _0202_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1145_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[105\] net109 _0691_
+ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1076_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[63\] net145 net128
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[79\] net98 vssd1 vssd1
+ vccd1 vccd1 _0657_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1673__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0929_ net270 _0018_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.nrst
+ sky130_fd_sc_hd__and2_2
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold13 net56 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[127\] vssd1 vssd1
+ vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[2\] vssd1 vssd1
+ vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net55 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold79 net57 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[126\] vssd1 vssd1
+ vccd1 vccd1 net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[118\] vssd1 vssd1
+ vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1832_ net236 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_38_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1763_ net190 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1694_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[9\]
+ net161 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout176_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1128_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[89\] net144 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[105\] net99 vssd1 vssd1
+ vccd1 vccd1 _0683_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1059_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[62\] net114 net89
+ _0648_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_36_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_12_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1815_ net154 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1746_ net241 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1677_ clknet_leaf_0_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[1\]
+ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input21_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1600_ clknet_leaf_22_wb_clk_i _0114_ net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1531_ clknet_leaf_24_wb_clk_i _0045_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1462_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[12\] _0346_ _0352_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[116\] _0384_ vssd1 vssd1
+ vccd1 vccd1 _0402_ sky130_fd_sc_hd__a221o_1
X_1393_ net118 net93 _0212_ _0322_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout139_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold110 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[98\] vssd1 vssd1
+ vccd1 vccd1 net370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1729_ clknet_leaf_12_wb_clk_i _0008_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold132 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[50\] vssd1 vssd1
+ vccd1 vccd1 net392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[20\] vssd1 vssd1
+ vccd1 vccd1 net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[39\] vssd1 vssd1
+ vccd1 vccd1 net381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0962_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[6\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[22\] vssd1 vssd1 vccd1
+ vccd1 _0600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0893_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[13\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__or4b_2
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1514_ clknet_leaf_14_wb_clk_i _0028_ net183 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1445_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[35\] _0342_ _0344_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[83\] vssd1 vssd1 vccd1
+ vccd1 _0386_ sky130_fd_sc_hd__a22o_1
X_1376_ _0209_ _0317_ _0318_ _0726_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout82 net84 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_2
XFILLER_0_36_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1834__237 vssd1 vssd1 vccd1 vccd1 _1834__237/HI net237 sky130_fd_sc_hd__conb_1
XFILLER_0_52_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1230_ team_11_WB.instance_to_wrap.sending.currentState\[5\] _0728_ _0214_ vssd1
+ vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__o21ba_2
Xclkbuf_leaf_26_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_1161_ net355 net109 net85 _0699_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__o22a_1
XANTENNA__1496__A2 _0346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1092_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[71\] net145 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[87\] net98 vssd1 vssd1
+ vccd1 vccd1 _0665_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0945_ net152 _0587_ _0460_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__o21ai_1
X_0876_ _0535_ _0540_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1428_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[33\] _0342_ _0349_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[17\] _0370_ vssd1 vssd1
+ vccd1 vccd1 _0371_ sky130_fd_sc_hd__a221o_1
XANTENNA__1596__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1359_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[13\] net152 net140
+ _0254_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0752__C net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1411__A2 _0345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1213_ team_11_WB.instance_to_wrap.sending.currentState\[0\] team_11_WB.instance_to_wrap.sending.currentState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1144_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[97\] net144 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[113\] net99 vssd1 vssd1
+ vccd1 vccd1 _0691_ sky130_fd_sc_hd__a221o_1
X_1075_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[70\] net114 net88
+ _0656_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout121_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0928_ team_11_WB.EN_VAL_REG net155 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__or2_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0859_ net296 _0527_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[26\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1783__206 vssd1 vssd1 vccd1 vccd1 _1783__206/HI net206 sky130_fd_sc_hd__conb_1
Xhold14 team_11_WB.instance_to_wrap.sending.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 team_11_WB.instance_to_wrap.sending.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net285 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold47 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[4\] vssd1 vssd1
+ vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[26\] vssd1 vssd1 vccd1 vccd1
+ net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[20\] vssd1 vssd1 vccd1 vccd1
+ net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[22\] vssd1 vssd1 vccd1 vccd1
+ net329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1831_ net153 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1762_ net189 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_53_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1693_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[8\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1771__198 vssd1 vssd1 vccd1 vccd1 _1771__198/HI net198 sky130_fd_sc_hd__conb_1
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1127_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[96\] net105 net83
+ _0682_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1058_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[54\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[70\] vssd1 vssd1 vccd1
+ vccd1 _0648_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1075__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1540__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1699__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1537__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1814_ net231 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_1745_ net240 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1676_ clknet_leaf_1_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[0\]
+ net157 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1789__212 vssd1 vssd1 vccd1 vccd1 _1789__212/HI net212 sky130_fd_sc_hd__conb_1
XANTENNA_input14_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1530_ clknet_leaf_14_wb_clk_i _0044_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_1461_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[100\] _0343_ _0349_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[20\] _0396_ vssd1 vssd1
+ vccd1 vccd1 _0401_ sky130_fd_sc_hd__a221o_1
X_1392_ net93 _0215_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__and3_4
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[68\] vssd1 vssd1
+ vccd1 vccd1 net360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1728_ clknet_leaf_12_wb_clk_i _0007_ net181 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold144 _0597_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[40\] vssd1 vssd1
+ vccd1 vccd1 net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[32\] vssd1 vssd1
+ vccd1 vccd1 net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 net48 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ clknet_leaf_7_wb_clk_i _0169_ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input6_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0961_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[13\] net105 net91
+ _0599_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1432__B1 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0892_ _0551_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1513_ clknet_leaf_2_wb_clk_i _0027_ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_1444_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[43\] _0336_ _0338_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[107\] vssd1 vssd1 vccd1
+ vccd1 _0385_ sky130_fd_sc_hd__a22o_1
X_1375_ net93 _0212_ _0321_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__and3_1
XANTENNA__1423__B1 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1827__234 vssd1 vssd1 vccd1 vccd1 _1827__234/HI net234 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_1_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout83 net84 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_2
XANTENNA__1414__B1 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout94 _0200_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1160_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[105\] net144 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[121\] vssd1 vssd1 vccd1
+ vccd1 _0699_ sky130_fd_sc_hd__a22o_1
XANTENNA_output45_A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[78\] net113 net88
+ _0664_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0944_ net152 _0587_ _0460_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0875_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[5\] _0539_ vssd1 vssd1 vccd1
+ vccd1 _0540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1184__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1427_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\] _0346_ _0352_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[113\] _0363_ vssd1 vssd1
+ vccd1 vccd1 _0370_ sky130_fd_sc_hd__a221o_1
X_1358_ net187 team_11_WB.instance_to_wrap.kp.controlstop.upper vssd1 vssd1 vccd1
+ vccd1 _0310_ sky130_fd_sc_hd__nand2_1
X_1289_ _0584_ _0240_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_26_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0998__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1212_ team_11_WB.instance_to_wrap.sending.currentState\[1\] net94 net135 vssd1 vssd1
+ vccd1 vccd1 _0145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1143_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[104\] net105 net83
+ _0690_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__o22a_1
X_1074_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[62\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[78\] vssd1 vssd1 vccd1
+ vccd1 _0656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1776__203 vssd1 vssd1 vccd1 vccd1 _1776__203/HI net203 sky130_fd_sc_hd__conb_1
XFILLER_0_62_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0927_ net388 _0576_ _0577_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0858_ _0526_ _0527_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[25\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0789_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[15\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold37 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[18\] vssd1 vssd1 vccd1 vccd1
+ net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 team_11_WB.instance_to_wrap.sending.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net275 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[0\] vssd1 vssd1
+ vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[11\] vssd1 vssd1 vccd1 vccd1
+ net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[124\] vssd1 vssd1
+ vccd1 vccd1 net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1148__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1830_ net235 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_53_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1761_ net256 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1692_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[7\]
+ net161 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_1126_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[88\] net140 net124
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[104\] vssd1 vssd1 vccd1
+ vccd1 _0682_ sky130_fd_sc_hd__a22o_1
X_1057_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[61\] net106 net91
+ _0647_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1813_ net154 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
X_1744_ net239 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1675_ clknet_leaf_24_wb_clk_i _0185_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout181_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1109_ net389 net104 _0673_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1460_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[52\] _0339_ _0347_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[28\] _0398_ vssd1 vssd1
+ vccd1 vccd1 _0400_ sky130_fd_sc_hd__a221o_1
X_1391_ net118 _0322_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold101 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[44\] vssd1 vssd1
+ vccd1 vccd1 net361 sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ clknet_leaf_12_wb_clk_i _0006_ net184 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold123 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[100\] vssd1 vssd1
+ vccd1 vccd1 net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 net45 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[59\] vssd1 vssd1
+ vccd1 vccd1 net372 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ clknet_leaf_7_wb_clk_i _0168_ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold145 _0026_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1589_ clknet_leaf_20_wb_clk_i _0103_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1804__224 vssd1 vssd1 vccd1 vccd1 _1804__224/HI net224 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0960_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[5\] net141 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[21\] vssd1 vssd1 vccd1
+ vccd1 _0599_ sky130_fd_sc_hd__a22o_1
XANTENNA__1432__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0891_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[9\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[11\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _0551_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1512_ clknet_leaf_23_wb_clk_i net405 net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_1443_ _0199_ _0214_ _0322_ _0557_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__a31o_1
X_1374_ _0213_ _0316_ _0322_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1187__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout95 net100 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_2
Xfanout84 net89 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_40_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1090_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[70\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[86\] vssd1 vssd1 vccd1
+ vccd1 _0664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0943_ team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl net140 vssd1 vssd1
+ vccd1 vccd1 _0587_ sky130_fd_sc_hd__or2_1
X_0874_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[4\] _0538_ vssd1 vssd1 vccd1
+ vccd1 _0539_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1426_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[121\] _0341_ _0348_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[73\] _0364_ vssd1 vssd1
+ vccd1 vccd1 _0369_ sky130_fd_sc_hd__a221o_1
X_1357_ _0441_ _0250_ _0255_ _0257_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__or4_1
X_1288_ _0238_ _0241_ _0244_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1753__248 vssd1 vssd1 vccd1 vccd1 net248 _1753__248/LO sky130_fd_sc_hd__conb_1
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1020__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1211_ _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__nand2_1
X_1142_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[96\] net140 net124
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[112\] vssd1 vssd1 vccd1
+ vccd1 _0690_ sky130_fd_sc_hd__a22o_1
X_1073_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[69\] net106 net91
+ _0655_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0926_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[14\] _0576_ _0558_ vssd1 vssd1
+ vccd1 vccd1 _0577_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0857_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[25\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[24\]
+ _0525_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__and3_1
X_0788_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[19\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[18\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[21\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout107_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold16 team_11_WB.instance_to_wrap.sending.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net276 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold27 _0150_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[104\] _0338_ _0343_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[96\] vssd1 vssd1 vccd1
+ vccd1 _0353_ sky130_fd_sc_hd__a22o_1
Xhold38 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[8\] vssd1 vssd1 vccd1 vccd1
+ net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[28\] vssd1 vssd1 vccd1 vccd1
+ net309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input37_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1760_ net255 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1691_ clknet_leaf_4_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[6\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1125_ net364 net104 _0681_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__o21a_1
X_1056_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[53\] net141 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[69\] vssd1 vssd1 vccd1
+ vccd1 _0647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0909_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\] _0563_ vssd1 vssd1 vccd1
+ vccd1 _0566_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1759__254 vssd1 vssd1 vccd1 vccd1 net254 _1759__254/LO sky130_fd_sc_hd__conb_1
XFILLER_0_54_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1462__C1 _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1812_ net153 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1743_ clknet_leaf_20_wb_clk_i _0002_ _0019_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
X_1674_ clknet_leaf_2_wb_clk_i _0184_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1108_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[79\] net138 net122
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[95\] net97 vssd1 vssd1
+ vccd1 vccd1 _0673_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1039_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[52\] net101 net82
+ _0638_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout87_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0970__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1390_ net56 _0328_ _0334_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_38_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1450__A2 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1726_ clknet_leaf_12_wb_clk_i _0005_ net184 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold102 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[79\] vssd1 vssd1
+ vccd1 vccd1 net362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[47\] vssd1 vssd1
+ vccd1 vccd1 net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[83\] vssd1 vssd1
+ vccd1 vccd1 net384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[72\] vssd1 vssd1
+ vccd1 vccd1 net395 sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ clknet_leaf_11_wb_clk_i _0167_ net181 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold146 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[54\] vssd1 vssd1
+ vccd1 vccd1 net406 sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ clknet_leaf_24_wb_clk_i _0102_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold134_A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0952__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0890_ _0541_ _0549_ _0550_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1432__A2 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1511_ clknet_leaf_17_wb_clk_i _0025_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1442_ net172 _0382_ _0383_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__and3_1
X_1373_ _0202_ _0203_ _0209_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_46_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1423__A2 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1709_ clknet_leaf_8_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[24\]
+ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_18_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_1_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_54_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1414__A2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout85 net89 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_2
Xfanout96 net100 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_2
XFILLER_0_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1767__194 vssd1 vssd1 vccd1 vccd1 _1767__194/HI net194 sky130_fd_sc_hd__conb_1
XANTENNA__1350__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0942_ team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl net136 vssd1 vssd1
+ vccd1 vccd1 _0586_ sky130_fd_sc_hd__nor2_1
X_0873_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[1\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[0\]
+ team_11_WB.instance_to_wrap.sending.cnt_20ms\[3\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1425_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[81\] _0344_ _0347_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[25\] _0365_ vssd1 vssd1
+ vccd1 vccd1 _0368_ sky130_fd_sc_hd__a221o_1
X_1356_ _0260_ _0276_ net90 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__a21oi_1
X_1287_ _0582_ _0216_ _0240_ _0714_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_46_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1574__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1210_ _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__and2_1
X_1141_ net385 net104 _0689_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1072_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[61\] net140 net124
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[77\] vssd1 vssd1 vccd1
+ vccd1 _0655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0925_ _0576_ _0541_ _0575_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__and3b_1
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0856_ net280 _0525_ net310 vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0787_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[27\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[26\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[29\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__or4_1
Xhold17 team_11_WB.instance_to_wrap.sending.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[14\] vssd1 vssd1 vccd1 vccd1
+ net288 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ _0199_ _0318_ _0321_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__and3_4
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold39 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[19\] vssd1 vssd1 vccd1 vccd1
+ net299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1339_ _0239_ _0292_ _0293_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1690_ clknet_leaf_4_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[5\]
+ net161 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1124_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[87\] net138 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[103\] net96 vssd1 vssd1
+ vccd1 vccd1 _0681_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1055_ net347 net101 _0646_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1480__B1 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0908_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\] _0563_ vssd1 vssd1 vccd1
+ vccd1 _0565_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0839_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[17\] _0484_ _0510_ vssd1 vssd1
+ vccd1 vccd1 _0517_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1471__B1 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1462__B1 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1811_ net153 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_13_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1742_ clknet_leaf_22_wb_clk_i _0198_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1673_ clknet_leaf_2_wb_clk_i _0183_ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1107_ net352 net114 net87 _0672_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_52_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1038_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[44\] net136 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[60\] vssd1 vssd1 vccd1
+ vccd1 _0638_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1796__219 vssd1 vssd1 vccd1 vccd1 _1796__219/HI net219 sky130_fd_sc_hd__conb_1
XFILLER_0_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1444__B1 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1435__B1 _0345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1725_ clknet_leaf_12_wb_clk_i _0004_ net184 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[33\] vssd1 vssd1
+ vccd1 vccd1 net363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold125 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[103\] vssd1 vssd1
+ vccd1 vccd1 net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[35\] vssd1 vssd1
+ vccd1 vccd1 net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 team_11_WB.instance_to_wrap.sending.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1
+ net407 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ clknet_leaf_7_wb_clk_i _0166_ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold136 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[73\] vssd1 vssd1
+ vccd1 vccd1 net396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1587_ clknet_leaf_23_wb_clk_i _0101_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1426__B1 _0348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1114__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1510_ clknet_leaf_19_wb_clk_i _0024_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1441_ net44 net135 vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1372_ net118 _0320_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__and2b_1
XANTENNA__1120__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1779__258 vssd1 vssd1 vccd1 vccd1 net258 _1779__258/LO sky130_fd_sc_hd__conb_1
XFILLER_0_46_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ clknet_leaf_3_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[23\]
+ net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_1639_ clknet_leaf_26_wb_clk_i team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl
+ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.controlstop.msg_tx_ctrl
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input4_A gpio_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1709__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout86 net89 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_2
Xfanout97 net100 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_40_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1810__230 vssd1 vssd1 vccd1 vccd1 _1810__230/HI net230 sky130_fd_sc_hd__conb_1
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0941_ _0458_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0872_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[1\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[0\]
+ team_11_WB.instance_to_wrap.sending.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _0537_
+ sky130_fd_sc_hd__and3_1
X_1424_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[1\] _0340_ _0343_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[97\] _0366_ vssd1 vssd1
+ vccd1 vccd1 _0367_ sky130_fd_sc_hd__a221o_1
X_1355_ net343 net90 _0306_ _0307_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__a22o_1
X_1286_ _0714_ _0240_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1140_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[95\] net137 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[111\] net100 vssd1 vssd1
+ vccd1 vccd1 _0689_ sky130_fd_sc_hd__a221o_1
X_1071_ net360 net101 _0654_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0924_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[13\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\]
+ _0572_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0855_ net280 _0525_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[24\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0786_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[23\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[22\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[25\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[24\]
+ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold29 team_11_WB.instance_to_wrap.sending.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 _0233_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ net118 net93 _0318_ _0322_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__and4_4
XTAP_TAPCELL_ROW_3_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1338_ _0242_ _0246_ net187 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__o21a_1
X_1269_ _0230_ _0231_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1724__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1123_ net365 net114 net87 _0680_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__o22a_1
X_1054_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[52\] net137 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[68\] net95 vssd1 vssd1
+ vccd1 vccd1 _0646_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0907_ net325 _0562_ _0564_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0838_ _0484_ _0510_ net334 vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__a21oi_1
X_0769_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[0\] team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1810_ net230 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_13_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1741_ clknet_leaf_14_wb_clk_i _0197_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1672_ clknet_leaf_25_wb_clk_i _0182_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1106_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[78\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[94\] vssd1 vssd1 vccd1
+ vccd1 _0672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1037_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[51\] net111 net87
+ _0637_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_52_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1724_ clknet_leaf_12_wb_clk_i _0017_ net184 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold104 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[95\] vssd1 vssd1
+ vccd1 vccd1 net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[31\] vssd1 vssd1
+ vccd1 vccd1 net375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[30\] vssd1 vssd1
+ vccd1 vccd1 net386 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ clknet_leaf_11_wb_clk_i _0165_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold148 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[13\] vssd1 vssd1 vccd1 vccd1
+ net408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold137 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[80\] vssd1 vssd1
+ vccd1 vccd1 net397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1586_ clknet_leaf_13_wb_clk_i _0100_ net183 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[86\]
+ sky130_fd_sc_hd__dfrtp_1
X_1749__244 vssd1 vssd1 vccd1 vccd1 net244 _1749__244/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_37_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1440_ _0375_ _0377_ _0379_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__or4_1
X_1371_ team_11_WB.instance_to_wrap.sending.currentState\[5\] _0208_ _0203_ _0202_
+ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1707_ clknet_leaf_8_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[22\]
+ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_1638_ clknet_leaf_15_wb_clk_i _0149_ net183 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.currentState\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_1569_ clknet_leaf_9_wb_clk_i _0083_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[69\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_1_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout98 net99 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_4
Xfanout87 net88 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_40_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0940_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[5\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[4\]
+ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[7\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__or4b_4
XFILLER_0_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0871_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[1\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1423_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[57\] _0350_ _0351_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[89\] vssd1 vssd1 vccd1
+ vccd1 _0366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1354_ _0261_ _0266_ net90 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__o21ba_1
X_1285_ _0582_ _0216_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_13_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout142_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1070_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[60\] net136 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[76\] net95 vssd1 vssd1
+ vccd1 vccd1 _0654_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0923_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\] _0572_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0854_ net291 _0524_ _0525_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[23\]
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0785_ net273 _0480_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold19 net54 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ _0215_ _0316_ _0322_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__and3_4
X_1337_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\] net152 _0257_
+ _0441_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1268_ net289 _0228_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__nor2_1
X_1199_ team_11_WB.instance_to_wrap.sending.currentState\[1\] team_11_WB.instance_to_wrap.sending.currentState\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1122_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[86\] net150 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[102\] vssd1 vssd1 vccd1
+ vccd1 _0680_ sky130_fd_sc_hd__a22o_1
X_1053_ net372 net113 _0645_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__o21a_1
XANTENNA__1628__SET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1480__A2 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0906_ _0535_ _0540_ _0563_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0837_ net330 _0513_ _0515_ _0491_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[16\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0768_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[5\] team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout105_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input35_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1462__A2 _0346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ clknet_leaf_15_wb_clk_i _0196_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1671_ clknet_leaf_24_wb_clk_i _0181_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1686__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1105_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[85\] net106 net92
+ _0671_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__o22a_1
X_1036_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[43\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[59\] vssd1 vssd1 vccd1
+ vccd1 _0637_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1444__A2 _0336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0955__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1435__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1723_ clknet_leaf_12_wb_clk_i _0016_ net184 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[25\] vssd1 vssd1
+ vccd1 vccd1 net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[94\] vssd1 vssd1
+ vccd1 vccd1 net365 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ clknet_leaf_11_wb_clk_i _0164_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold138 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[65\] vssd1 vssd1
+ vccd1 vccd1 net398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold127 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[114\] vssd1 vssd1
+ vccd1 vccd1 net387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[1\] vssd1 vssd1 vccd1 vccd1
+ net409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1585_ clknet_leaf_9_wb_clk_i _0099_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[85\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout172_A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1426__A2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1019_ net366 net111 _0628_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout85_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1370_ _0209_ _0317_ _0318_ _0557_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1706_ clknet_leaf_6_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[21\]
+ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_1637_ clknet_leaf_10_wb_clk_i _0148_ net178 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.currentState\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_1786__209 vssd1 vssd1 vccd1 vccd1 _1786__209/HI net209 sky130_fd_sc_hd__conb_1
X_1568_ clknet_leaf_22_wb_clk_i _0082_ net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1499_ _0428_ _0430_ _0433_ _0435_ net170 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__o41ai_1
XTAP_TAPCELL_ROW_1_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout99 net100 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_4
Xfanout88 net89 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_2
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0870_ _0532_ _0533_ _0534_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1422_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[49\] _0339_ _0345_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[65\] vssd1 vssd1 vccd1
+ vccd1 _0365_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_50_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1353_ _0249_ _0253_ _0277_ _0305_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a31o_1
X_1284_ _0714_ _0216_ _0240_ _0582_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__o22ai_2
XTAP_TAPCELL_ROW_47_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout135_A _0556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0999_ net393 net115 net88 _0618_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1813__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1552__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1492__B1 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0922_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\] _0572_ _0574_ vssd1 vssd1
+ vccd1 vccd1 _0006_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0853_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[21\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[23\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[22\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0525_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0784_ net284 _0480_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[2\]
+ sky130_fd_sc_hd__nor2_1
X_1405_ net94 _0215_ _0321_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__and3_4
X_1336_ _0264_ _0289_ _0291_ _0275_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__a31o_1
Xinput1 gpio_in[34] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
X_1267_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[12\] _0228_ vssd1 vssd1 vccd1
+ vccd1 _0230_ sky130_fd_sc_hd__and2_1
X_1198_ team_11_WB.instance_to_wrap.sending.currentState\[1\] _0439_ _0440_ _0716_
+ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__1483__B1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1474__B1 _0348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1561__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1121_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[93\] net105 net91
+ _0679_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__o22a_1
X_1052_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[51\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[67\] net98 vssd1 vssd1
+ vccd1 vccd1 _0645_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0905_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[7\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[6\]
+ _0559_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0836_ _0484_ _0510_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1830__235 vssd1 vssd1 vccd1 vccd1 _1830__235/HI net235 sky130_fd_sc_hd__conb_1
X_0767_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[6\] team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1319_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[1\] net90 vssd1 vssd1
+ vccd1 vccd1 _0275_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1456__B1 _0342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1144__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1447__B1 _0349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1212__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1670_ clknet_leaf_24_wb_clk_i _0180_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1104_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[77\] net143 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[93\] vssd1 vssd1 vccd1
+ vccd1 _0671_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1035_ net392 net111 net86 _0636_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__o22a_1
XANTENNA__1438__B1 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0819_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[10\] _0498_ _0501_ vssd1 vssd1
+ vccd1 vccd1 _0504_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1799_ net222 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XANTENNA__1821__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1132__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1722_ clknet_leaf_11_wb_clk_i _0015_ net181 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1653_ clknet_leaf_11_wb_clk_i _0163_ net181 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold106 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[42\] vssd1 vssd1
+ vccd1 vccd1 net366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[71\] vssd1 vssd1
+ vccd1 vccd1 net377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold128 team_11_WB.instance_to_wrap.sending.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1
+ net388 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold139 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[92\] vssd1 vssd1
+ vccd1 vccd1 net399 sky130_fd_sc_hd__dlygate4sd3_1
X_1584_ clknet_leaf_22_wb_clk_i _0098_ net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout165_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1018_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[34\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[50\] net99 vssd1 vssd1
+ vccd1 vccd1 _0628_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1816__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1506__RESET_B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1180__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1705_ clknet_leaf_6_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[20\]
+ net166 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1755__250 vssd1 vssd1 vccd1 vccd1 net250 _1755__250/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_57_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1636_ clknet_leaf_10_wb_clk_i _0147_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.currentState\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_1567_ clknet_leaf_18_wb_clk_i _0081_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_1498_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[95\] _0351_ _0426_
+ _0427_ _0434_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__a2111o_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout89 _0592_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1421_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[41\] _0336_ _0338_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[105\] vssd1 vssd1 vccd1
+ vccd1 _0364_ sky130_fd_sc_hd__a22o_1
X_1352_ net188 _0251_ _0252_ _0284_ _0304_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a311o_1
X_1283_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[0\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[2\]
+ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[3\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_47_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout128_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0998_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[24\] net150 net133
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[40\] vssd1 vssd1 vccd1
+ vccd1 _0618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1619_ clknet_leaf_23_wb_clk_i _0133_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input2_A gpio_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1521__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0921_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\] _0572_ _0541_ vssd1 vssd1
+ vccd1 vccd1 _0574_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0852_ _0523_ _0524_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[22\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0783_ net279 _0480_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1404_ _0199_ _0318_ _0335_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__and3_4
X_1335_ _0261_ _0281_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__or2_1
Xinput2 gpio_in[35] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_1
X_1266_ _0228_ _0229_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1197_ team_11_WB.instance_to_wrap.sending.currentState\[1\] team_11_WB.instance_to_wrap.sending.currentState\[2\]
+ team_11_WB.instance_to_wrap.sending.currentState\[0\] vssd1 vssd1 vccd1 vccd1 _0719_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__1483__B2 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1171__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1702__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1120_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[85\] net143 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[101\] vssd1 vssd1 vccd1
+ vccd1 _0679_ sky130_fd_sc_hd__a22o_1
X_1051_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[58\] net111 net86
+ _0644_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0904_ _0562_ net117 _0561_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0835_ _0491_ _0512_ _0514_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[15\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_43_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0766_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[1\] team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1318_ net90 _0272_ _0274_ _0265_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__o31a_1
X_1249_ _0538_ _0220_ net117 vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__o21bai_1
X_1763__190 vssd1 vssd1 vccd1 vccd1 _1763__190/HI net190 sky130_fd_sc_hd__conb_1
XFILLER_0_63_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1819__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1807__227 vssd1 vssd1 vccd1 vccd1 _1807__227/HI net227 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_54_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1080__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1103_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[84\] net101 net82
+ _0670_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__o22a_1
X_1034_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[42\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[58\] vssd1 vssd1 vccd1
+ vccd1 _0636_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1798_ net221 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
X_0818_ _0491_ _0500_ _0503_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[9\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0749_ net30 net29 _0452_ _0453_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input40_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1721_ clknet_leaf_11_wb_clk_i _0014_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1652_ clknet_leaf_11_wb_clk_i _0162_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold107 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[107\] vssd1 vssd1
+ vccd1 vccd1 net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[28\] vssd1 vssd1
+ vccd1 vccd1 net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[87\] vssd1 vssd1
+ vccd1 vccd1 net389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1583_ clknet_leaf_18_wb_clk_i _0097_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1017_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[41\] net109 net84
+ _0627_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout158_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1704_ clknet_leaf_6_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[19\]
+ net166 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1635_ clknet_leaf_10_wb_clk_i _0146_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.currentState\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1566_ clknet_leaf_20_wb_clk_i _0080_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1497_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[31\] _0347_ _0349_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[23\] vssd1 vssd1 vccd1
+ vccd1 _0434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1727__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1420_ net118 net93 _0212_ _0320_ _0557_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__a41o_1
X_1351_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[12\] _0583_ _0245_
+ _0441_ _0258_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__a221o_1
X_1282_ _0714_ _0216_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1792__215 vssd1 vssd1 vccd1 vccd1 _1792__215/HI net215 sky130_fd_sc_hd__conb_1
XFILLER_0_61_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0997_ net375 net101 _0617_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1618_ clknet_leaf_15_wb_clk_i _0132_ net183 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1549_ clknet_leaf_21_wb_clk_i _0063_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1492__A2 _0336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1231__S _0556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0920_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[11\] _0569_ _0573_ _0558_ vssd1
+ vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__o211a_1
X_0851_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[21\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[22\]
+ _0522_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0782_ net321 _0480_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1403_ net118 net93 _0215_ _0320_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__and4_4
X_1334_ _0249_ _0260_ net90 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__a21oi_1
X_1265_ net407 _0226_ net276 vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__a21oi_1
Xinput3 gpio_in[36] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
X_1196_ team_11_WB.instance_to_wrap.sending.currentState\[2\] _0717_ vssd1 vssd1 vccd1
+ vccd1 _0718_ sky130_fd_sc_hd__xnor2_1
XANTENNA__1483__A2 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout140_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1474__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1050_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[50\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[66\] vssd1 vssd1 vccd1
+ vccd1 _0644_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1465__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0903_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[6\] _0559_ vssd1 vssd1 vccd1
+ vccd1 _0562_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0834_ _0513_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0765_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[7\] team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_47_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1317_ _0257_ _0266_ _0268_ _0273_ _0591_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a2111o_1
X_1248_ net320 _0537_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1456__A2 _0336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1798__221 vssd1 vssd1 vccd1 vccd1 _1798__221/HI net221 sky130_fd_sc_hd__conb_1
XFILLER_0_63_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1179_ net305 net112 net86 _0708_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1835__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1447__A2 _0345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1102_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[76\] net137 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[92\] vssd1 vssd1 vccd1
+ vccd1 _0670_ sky130_fd_sc_hd__a22o_1
X_1033_ net358 net103 net84 _0635_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1438__A2 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1797_ net220 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0817_ _0502_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__inv_2
X_0748_ net26 net27 vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout103_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input33_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1720_ clknet_leaf_12_wb_clk_i _0013_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1651_ clknet_leaf_11_wb_clk_i _0161_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold108 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[48\] vssd1 vssd1
+ vccd1 vccd1 net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[57\] vssd1 vssd1
+ vccd1 vccd1 net379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1582_ clknet_leaf_19_wb_clk_i _0096_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1016_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[33\] net144 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[49\] vssd1 vssd1 vccd1
+ vccd1 _0627_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_16_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1347__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1515__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1703_ clknet_leaf_6_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[18\]
+ net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1634_ clknet_leaf_13_wb_clk_i _0145_ net183 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.currentState\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1565_ clknet_leaf_21_wb_clk_i _0079_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_1496_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[15\] _0346_ _0431_
+ _0432_ _0326_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout170_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1017__B1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout83_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1350_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[3\] net90 _0290_
+ _0303_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__a22o_1
X_1281_ _0714_ _0237_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__nor2_1
XANTENNA__1495__B1 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0996_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[23\] net138 net120
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[39\] net96 vssd1 vssd1
+ vccd1 vccd1 _0617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1617_ clknet_leaf_10_wb_clk_i _0131_ net178 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[117\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1548_ clknet_leaf_15_wb_clk_i _0062_ net178 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_1479_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[78\] _0348_ _0349_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[22\] vssd1 vssd1 vccd1
+ vccd1 _0417_ sky130_fd_sc_hd__a22o_1
XANTENNA__1486__B1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1838__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1410__B1 _0348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1745__240 vssd1 vssd1 vccd1 vccd1 net240 _1745__240/LO sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0850_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[21\] _0522_ net329 vssd1 vssd1
+ vccd1 vccd1 _0523_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0781_ _0480_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keyvalid
+ sky130_fd_sc_hd__inv_2
XFILLER_0_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1402_ _0199_ _0215_ _0321_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__and3_4
X_1333_ _0286_ _0287_ _0288_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__or3_1
X_1264_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[10\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[11\]
+ _0226_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__and3_1
Xinput4 gpio_in[37] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_1
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1468__B1 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1195_ team_11_WB.instance_to_wrap.sending.currentState\[3\] team_11_WB.instance_to_wrap.sending.currentState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout133_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0979_ net354 net113 net87 _0608_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1459__B1 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1711__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0902_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[6\] _0559_ vssd1 vssd1 vccd1
+ vccd1 _0561_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0833_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[15\] _0510_ vssd1 vssd1 vccd1
+ vccd1 _0513_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0764_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[3\] team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1316_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[8\] net152 _0249_
+ _0255_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__a22o_1
X_1247_ _0537_ _0219_ net117 vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1178_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[114\] net147 vssd1
+ vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1101_ net384 net113 _0669_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__o21a_1
X_1032_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[41\] net137 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[57\] vssd1 vssd1 vccd1
+ vccd1 _0635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
X_1796_ net219 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0816_ _0498_ _0501_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__and2_1
XANTENNA__1633__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0747_ net23 net22 net25 net24 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input26_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1650_ clknet_leaf_11_wb_clk_i _0160_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1581_ clknet_leaf_21_wb_clk_i _0095_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[81\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold109 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[26\] vssd1 vssd1
+ vccd1 vccd1 net369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1015_ net371 net107 net84 _0626_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1779_ net258 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_13_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1702_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[17\]
+ net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1633_ clknet_leaf_13_wb_clk_i _0144_ net184 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.currentState\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1564_ clknet_leaf_16_wb_clk_i _0078_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_1495_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[79\] _0348_ _0352_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[119\] vssd1 vssd1 vccd1
+ vccd1 _0432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout163_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1280_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[1\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[2\]
+ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[3\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__or4b_4
XFILLER_0_25_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0995_ net386 net113 net87 _0616_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1616_ clknet_leaf_23_wb_clk_i _0130_ net169 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1547_ clknet_leaf_16_wb_clk_i _0061_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_1478_ _0410_ _0415_ _0416_ net178 vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0780_ net2 net1 net4 net3 vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nor4_2
XFILLER_0_24_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1401_ _0316_ _0318_ _0322_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__and3_4
XANTENNA__1165__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1332_ _0253_ _0282_ _0283_ _0285_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a211o_1
X_1263_ net281 _0226_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__xor2_1
Xinput5 wb_rst_i vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_1
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1194_ team_11_WB.instance_to_wrap.sending.currentState\[3\] team_11_WB.instance_to_wrap.sending.currentState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0978_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[30\] vssd1 vssd1 vccd1
+ vccd1 _0608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1782__205 vssd1 vssd1 vccd1 vccd1 _1782__205/HI net205 sky130_fd_sc_hd__conb_1
XFILLER_0_56_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0901_ _0559_ _0560_ _0558_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0832_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[15\] _0510_ vssd1 vssd1 vccd1
+ vccd1 _0512_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0763_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[4\] team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1315_ _0252_ _0269_ _0270_ _0271_ net187 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__o41a_1
X_1246_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[1\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[0\]
+ net327 vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a21oi_1
X_1177_ net313 net109 net85 _0707_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1770__197 vssd1 vssd1 vccd1 vccd1 _1770__197/HI net197 sky130_fd_sc_hd__conb_1
XFILLER_0_30_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1509__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1781__260 vssd1 vssd1 vccd1 vccd1 net260 _1781__260/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_54_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1100_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[75\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[91\] net98 vssd1 vssd1
+ vccd1 vccd1 _0669_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1031_ net368 net107 net84 _0634_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1639__D team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
X_1795_ net218 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_52_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput41 wbs_we_i vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0815_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[7\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[8\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[9\] vssd1 vssd1 vccd1 vccd1 _0501_
+ sky130_fd_sc_hd__and3_1
X_0746_ net15 net16 net13 net14 vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1229_ _0716_ _0205_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input19_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1580_ clknet_leaf_9_wb_clk_i _0094_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_1788__211 vssd1 vssd1 vccd1 vccd1 _1788__211/HI net211 sky130_fd_sc_hd__conb_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1491__B _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1014_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[32\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[48\] vssd1 vssd1 vccd1
+ vccd1 _0626_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_14_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1778_ net257 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1701_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[16\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1632_ clknet_leaf_1_wb_clk_i net263 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.debouncertop.next_receive_ready
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1563_ clknet_leaf_17_wb_clk_i _0077_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1494_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[55\] _0339_ _0345_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[71\] vssd1 vssd1 vccd1
+ vccd1 _0431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1705__RESET_B net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1495__A2 _0348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0994_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[22\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[38\] vssd1 vssd1 vccd1
+ vccd1 _0616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1615_ clknet_leaf_16_wb_clk_i _0129_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1546_ clknet_leaf_14_wb_clk_i _0060_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1477_ net47 _0556_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__or2_1
XANTENNA__1486__A2 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1410__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1400_ net93 _0318_ _0335_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__and3_4
X_1331_ _0249_ _0252_ _0276_ _0243_ _0280_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__a221o_1
X_1262_ _0226_ _0227_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__and2b_1
Xinput6 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA__1468__A2 _0342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1193_ net262 team_11_WB.instance_to_wrap.kp.debouncertop.receive_ready net157 vssd1
+ vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1698__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0977_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[21\] net106 net91
+ _0607_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout119_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1529_ clknet_leaf_9_wb_clk_i _0043_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[29\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1459__A2 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1775__202 vssd1 vssd1 vccd1 vccd1 _1775__202/HI net202 sky130_fd_sc_hd__conb_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0928__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[4\] _0547_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0831_ _0510_ _0511_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0762_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[2\] team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1314_ _0238_ _0241_ _0267_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__o21a_1
X_1245_ _0536_ _0218_ net117 vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__a21o_1
X_1176_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[113\] net145 vssd1
+ vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0930__C net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1030_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[40\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[56\] vssd1 vssd1 vccd1
+ vccd1 _0634_ sky130_fd_sc_hd__a22o_1
XANTENNA__1489__B _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput31 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0814_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[7\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[8\]
+ _0498_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _0500_ sky130_fd_sc_hd__a31o_1
X_1794_ net217 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0745_ net19 net18 net21 net20 vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1228_ team_11_WB.instance_to_wrap.sending.currentState\[4\] _0213_ net135 vssd1
+ vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1159_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[112\] net105 net83
+ _0698_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout99_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1013_ net381 net104 _0625_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_1_0__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1777_ net204 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout101_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input31_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1431__B1 _0348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1700_ clknet_leaf_5_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[15\]
+ net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1631_ clknet_leaf_25_wb_clk_i _0142_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.controlstop.mode
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1562_ clknet_leaf_14_wb_clk_i _0076_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1493_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[7\] _0340_ _0344_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[87\] _0429_ vssd1 vssd1
+ vccd1 vccd1 _0430_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1422__B1 _0345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1829_ net153 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1413__B1 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0993_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[29\] net106 net91
+ _0615_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1614_ clknet_leaf_18_wb_clk_i _0128_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1545_ clknet_leaf_8_wb_clk_i _0059_ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[45\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1476_ _0407_ _0411_ _0414_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1752__247 vssd1 vssd1 vccd1 vccd1 net247 _1752__247/LO sky130_fd_sc_hd__conb_1
XFILLER_0_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1330_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\] net152 _0279_
+ _0284_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__a211o_1
X_1261_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[7\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[8\]
+ _0223_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ _0227_ sky130_fd_sc_hd__a31o_1
Xinput7 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_1192_ _0441_ _0715_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0976_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[13\] net141 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[29\] vssd1 vssd1 vccd1
+ vccd1 _0607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1528_ clknet_leaf_23_wb_clk_i _0042_ net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_1459_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[108\] _0338_ _0340_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[4\] _0397_ vssd1 vssd1
+ vccd1 vccd1 _0399_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0830_ net408 _0508_ net288 vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0761_ _0462_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1313_ _0020_ _0246_ _0248_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__and3_1
X_1244_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[1\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__or2_1
X_1175_ net322 net105 net83 _0706_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0959_ team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl _0590_ net96 vssd1
+ vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1758__253 vssd1 vssd1 vccd1 vccd1 net253 _1758__253/LO sky130_fd_sc_hd__conb_1
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput10 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0813_ net298 _0499_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[8\]
+ sky130_fd_sc_hd__xnor2_1
X_1793_ net216 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0744_ _0445_ _0446_ _0447_ _0448_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1227_ _0212_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout179_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1158_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[104\] net140 net124
+ net322 vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1089_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[77\] net105 net92
+ _0663_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1611__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1012_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[31\] net138 net122
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[47\] net97 vssd1 vssd1
+ vccd1 vccd1 _0625_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1776_ net203 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input24_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1630_ clknet_leaf_3_wb_clk_i net261 net157 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.debouncertop.receive_ready
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1561_ clknet_leaf_9_wb_clk_i _0075_ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[61\]
+ sky130_fd_sc_hd__dfstp_1
X_1492_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[47\] _0336_ _0338_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[111\] vssd1 vssd1 vccd1
+ vccd1 _0429_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1828_ net154 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_20_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1759_ net254 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_40_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1714__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0992_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[21\] net140 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[37\] vssd1 vssd1 vccd1
+ vccd1 _0615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1613_ clknet_leaf_21_wb_clk_i _0127_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1544_ clknet_leaf_26_wb_clk_i _0058_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_1475_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[93\] _0351_ _0412_
+ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__a211o_1
X_1766__193 vssd1 vssd1 vccd1 vccd1 _1766__193/HI net193 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_25_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout161_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1260_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[7\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[9\]
+ team_11_WB.instance_to_wrap.sending.cnt_20ms\[8\] _0223_ vssd1 vssd1 vccd1 vccd1
+ _0226_ sky130_fd_sc_hd__and4_1
Xinput8 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
X_1191_ _0458_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0975_ net356 net101 net82 _0606_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1527_ clknet_leaf_18_wb_clk_i _0041_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_1458_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[68\] _0345_ _0348_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[76\] vssd1 vssd1 vccd1
+ vccd1 _0398_ sky130_fd_sc_hd__a22o_1
X_1389_ net55 _0329_ net53 net54 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1068__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0760_ team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[3\] net186
+ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
X_1312_ _0001_ _0021_ _0253_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__o21a_1
X_1243_ _0535_ _0540_ net274 vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1174_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[112\] net140 vssd1
+ vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0958_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[12\] net102 net82
+ net404 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout124_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0889_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[4\] _0547_ vssd1 vssd1 vccd1
+ vccd1 _0550_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1558__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput11 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0812_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[7\] _0498_ _0499_ _0491_ vssd1
+ vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[7\] sky130_fd_sc_hd__o211a_1
X_1792_ net215 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0743_ net10 net9 net12 net11 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1226_ _0440_ _0207_ _0211_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__o21ai_4
X_1157_ net390 net102 _0697_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1088_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[69\] net141 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[85\] vssd1 vssd1 vccd1
+ vccd1 _0663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_1011_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[38\] net113 net87
+ _0624_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_37_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1795__218 vssd1 vssd1 vccd1 vccd1 _1795__218/HI net218 sky130_fd_sc_hd__conb_1
XFILLER_0_60_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1775_ net202 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1209_ team_11_WB.instance_to_wrap.sending.currentState\[0\] _0718_ _0728_ team_11_WB.instance_to_wrap.sending.currentState\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input17_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1431__A2 _0336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1560_ clknet_leaf_22_wb_clk_i _0074_ net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1491_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[63\] _0350_ vssd1
+ vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1498__A2 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1422__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1827_ net234 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_5_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1758_ net253 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_1689_ clknet_leaf_4_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[4\]
+ net161 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input9_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1778__257 vssd1 vssd1 vccd1 vccd1 net257 _1778__257/LO sky130_fd_sc_hd__conb_1
XFILLER_0_36_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1413__A2 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0991_ net378 net101 _0614_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1612_ clknet_leaf_24_wb_clk_i _0126_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1543_ clknet_leaf_18_wb_clk_i _0057_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1474_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[53\] _0339_ _0348_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[77\] vssd1 vssd1 vccd1
+ vccd1 _0413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1190_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[4\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[6\]
+ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[7\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__or4b_4
Xinput9 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA_output48_A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0974_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[12\] net136 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[28\] vssd1 vssd1 vccd1
+ vccd1 _0606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1526_ clknet_leaf_21_wb_clk_i _0040_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1457_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[60\] _0350_ _0351_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[92\] vssd1 vssd1 vccd1
+ vccd1 _0397_ sky130_fd_sc_hd__a22o_1
X_1388_ net55 _0328_ _0333_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1311_ net187 _0267_ _0244_ _0260_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1242_ net265 _0217_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1173_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[119\] net102 _0705_
+ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1059__B1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0957_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[4\] net136 net119
+ net403 vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0888_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[4\] _0547_ vssd1 vssd1 vccd1
+ vccd1 _0549_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1545__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1509_ clknet_leaf_23_wb_clk_i _0023_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_54_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1470__B1 _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1598__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1461__B1 _0349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1791_ net214 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
Xinput12 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0811_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[7\] _0498_ vssd1 vssd1 vccd1
+ vccd1 _0499_ sky130_fd_sc_hd__nand2_1
Xinput34 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
X_0742_ net37 net36 net8 net7 vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or4_1
Xinput23 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1225_ team_11_WB.instance_to_wrap.sending.currentState\[3\] _0439_ _0728_ team_11_WB.instance_to_wrap.sending.currentState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a31o_1
X_1156_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[103\] net138 net120
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[119\] net96 vssd1 vssd1
+ vccd1 vccd1 _0697_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1087_ net342 net101 _0662_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1452__B1 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1691__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1140__C1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1708__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1010_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[30\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[46\] vssd1 vssd1 vccd1
+ vccd1 _0624_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1434__B1 _0349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1774_ net201 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout184_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1208_ team_11_WB.instance_to_wrap.sending.currentState\[0\] team_11_WB.instance_to_wrap.sending.currentState\[2\]
+ _0440_ _0716_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a2111o_1
X_1139_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[102\] net114 net87
+ _0688_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1425__B1 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout97_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1748__243 vssd1 vssd1 vccd1 vccd1 net243 _1748__243/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1416__B1 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1490_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[39\] _0342_ _0343_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[103\] vssd1 vssd1 vccd1
+ vccd1 _0427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1 team_11_WB.instance_to_wrap.kp.debouncertop.keyvalid vssd1 vssd1 vccd1 vccd1
+ net261 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1826_ net154 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1757_ net252 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1688_ clknet_leaf_4_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[3\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0990_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[20\] net136 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[36\] net95 vssd1 vssd1
+ vccd1 vccd1 _0614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1723__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1611_ clknet_leaf_23_wb_clk_i _0125_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1542_ clknet_leaf_20_wb_clk_i _0056_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1473_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[125\] _0341_ _0345_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[69\] vssd1 vssd1 vccd1
+ vccd1 _0412_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1809_ net229 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0973_ net344 net109 _0605_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1525_ clknet_leaf_23_wb_clk_i _0039_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_1456_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[44\] _0336_ _0342_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[36\] vssd1 vssd1 vccd1
+ vccd1 _0396_ sky130_fd_sc_hd__a22o_1
X_1387_ net54 _0330_ net53 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_18_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1310_ _0020_ _0248_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1241_ _0457_ _0216_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1172_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[111\] net139 net120
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[127\] net96 vssd1 vssd1
+ vccd1 vccd1 _0705_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0956_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\] net110 net85
+ _0596_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__o22a_1
X_0887_ net117 _0546_ _0548_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1508_ clknet_leaf_24_wb_clk_i _0022_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1439_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[98\] _0343_ _0350_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[58\] _0380_ vssd1 vssd1
+ vccd1 vccd1 _0381_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_54_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1790_ net213 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_52_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0810_ net269 _0496_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[6\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0741_ net17 net6 net31 net28 vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__or4_1
Xinput35 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
Xinput24 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1224_ team_11_WB.instance_to_wrap.sending.currentState\[3\] _0209_ net135 vssd1
+ vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__mux2_1
X_1155_ net357 net114 net87 _0696_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__o22a_1
X_1086_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[68\] net136 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[84\] net95 vssd1 vssd1
+ vccd1 vccd1 _0662_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0939_ _0458_ _0582_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0963__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1434__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1773_ net200 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1207_ team_11_WB.instance_to_wrap.sending.currentState\[0\] team_11_WB.instance_to_wrap.sending.currentState\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout177_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1138_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[94\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[110\] vssd1 vssd1 vccd1
+ vccd1 _0688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1069_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[67\] net113 _0653_
+ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1582__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold2 team_11_WB.instance_to_wrap.kp.debouncertop.next_receive_ready vssd1 vssd1
+ vccd1 vccd1 net262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1825_ net153 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1756_ net251 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1687_ clknet_leaf_3_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[2\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1785__208 vssd1 vssd1 vccd1 vccd1 _1785__208/HI net208 sky130_fd_sc_hd__conb_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input22_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1098__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1610_ clknet_leaf_13_wb_clk_i _0124_ net183 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1541_ clknet_leaf_21_wb_clk_i _0055_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1472_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[109\] _0338_ _0350_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[61\] _0406_ vssd1 vssd1
+ vccd1 vccd1 _0411_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1808_ net228 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_26_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1739_ clknet_leaf_22_wb_clk_i _0195_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0972_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\] net145 net128
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[27\] net98 vssd1 vssd1
+ vccd1 vccd1 _0605_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1524_ clknet_leaf_16_wb_clk_i _0038_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_1455_ net394 net135 net174 _0395_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__o211a_1
X_1386_ net53 _0331_ _0332_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1240_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[1\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[0\]
+ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[3\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__or4b_4
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1171_ net328 net115 net88 _0704_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0955_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[3\] net145 net128
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[19\] vssd1 vssd1 vccd1
+ vccd1 _0596_ sky130_fd_sc_hd__a22o_1
X_0886_ _0444_ _0545_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1507_ clknet_leaf_27_wb_clk_i _0021_ net160 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1438_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[82\] _0344_ _0352_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[114\] vssd1 vssd1 vccd1
+ vccd1 _0380_ sky130_fd_sc_hd__a22o_1
X_1369_ _0212_ _0215_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_54_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1470__A2 _0346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1536__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1461__A2 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput36 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
X_0740_ net33 net32 net35 net34 vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__or4_1
Xinput14 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0972__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1223_ team_11_WB.instance_to_wrap.sending.currentState\[5\] _0208_ vssd1 vssd1 vccd1
+ vccd1 _0210_ sky130_fd_sc_hd__or2_1
X_1154_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[102\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[118\] vssd1 vssd1 vccd1
+ vccd1 _0696_ sky130_fd_sc_hd__a22o_1
X_1085_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[75\] net113 _0661_
+ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout122_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0938_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[5\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[6\]
+ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[7\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__or4b_4
XFILLER_0_30_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0869_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[7\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[6\]
+ team_11_WB.instance_to_wrap.sending.cnt_20ms\[9\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0963__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0954__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1434__A2 _0346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1772_ net199 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1206_ _0727_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__inv_2
X_1137_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[101\] net108 net91
+ _0687_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1068_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[59\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[75\] net99 vssd1 vssd1
+ vccd1 vccd1 _0653_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1425__A2 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1416__A2 _0346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold3 _0143_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1824_ net233 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1755_ net250 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1686_ clknet_leaf_3_wb_clk_i net316 net163 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1639__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1031__B1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1540_ clknet_leaf_16_wb_clk_i _0054_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1471_ _0212_ _0317_ _0352_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[117\]
+ _0409_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1807_ net227 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1738_ clknet_leaf_18_wb_clk_i _0194_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1669_ clknet_leaf_25_wb_clk_i _0179_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ net331 net110 net85 _0604_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1523_ clknet_leaf_24_wb_clk_i _0037_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_1454_ _0386_ _0388_ _0391_ _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__or4_1
X_1385_ net54 _0328_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__or2_1
XANTENNA__1482__B1 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1473__B1 _0345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1170_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[110\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[126\] vssd1 vssd1 vccd1
+ vccd1 _0704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1839__238 vssd1 vssd1 vccd1 vccd1 _1839__238/HI net238 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_15_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0954_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\] net110 net85
+ _0595_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__o22a_1
X_0885_ _0444_ _0545_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1506_ clknet_leaf_27_wb_clk_i _0020_ net160 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1437_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[106\] _0338_ _0342_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[34\] _0378_ vssd1 vssd1
+ vccd1 vccd1 _0379_ sky130_fd_sc_hd__a221o_1
X_1368_ net118 _0729_ _0730_ _0204_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__and4_2
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1299_ _0584_ _0216_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1446__B1 _0348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput37 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xinput26 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1222_ team_11_WB.instance_to_wrap.sending.currentState\[3\] _0205_ _0206_ _0440_
+ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__o211a_2
X_1806__226 vssd1 vssd1 vccd1 vccd1 _1806__226/HI net226 sky130_fd_sc_hd__conb_1
X_1153_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[109\] net107 net92
+ _0695_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__o22a_1
X_1084_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[67\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[83\] net98 vssd1 vssd1
+ vccd1 vccd1 _0661_ sky130_fd_sc_hd__a221o_1
XANTENNA__1437__B1 _0342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0937_ _0581_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0868_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[13\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[12\]
+ team_11_WB.instance_to_wrap.sending.cnt_20ms\[10\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_30_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0799_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[1\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[0\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[2\] vssd1 vssd1 vccd1 vccd1 _0492_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1428__B1 _0349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout181 net185 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1840_ net153 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1771_ net198 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1205_ _0437_ _0724_ net135 vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1122__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1136_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[93\] net143 net126
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[109\] vssd1 vssd1 vccd1
+ vccd1 _0687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1067_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[66\] net111 net86
+ _0652_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_21_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 team_11_WB.instance_to_wrap.sending.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net264 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1104__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1591__RESET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1520__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1823_ net154 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1754_ net249 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1685_ clknet_leaf_3_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[0\]
+ net161 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1119_ net399 net103 net82 _0678_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout95_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1470_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[13\] _0346_ _0384_
+ _0405_ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1701__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1806_ net226 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1737_ clknet_leaf_20_wb_clk_i _0193_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1668_ clknet_leaf_2_wb_clk_i _0178_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1599_ clknet_leaf_17_wb_clk_i _0113_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_37_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1791__214 vssd1 vssd1 vccd1 vccd1 _1791__214/HI net214 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1205__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0970_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\] net147 net128
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[26\] vssd1 vssd1 vccd1
+ vccd1 _0604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1522_ clknet_leaf_14_wb_clk_i _0036_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_1453_ _0324_ _0385_ _0392_ _0393_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__or4_1
X_1384_ _0328_ _0331_ net53 vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout145_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0953_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[2\] net147 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[18\] vssd1 vssd1 vccd1
+ vccd1 _0595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0884_ _0444_ _0545_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1505_ net5 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1436_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[26\] _0347_ _0351_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[90\] vssd1 vssd1 vccd1
+ vccd1 _0378_ sky130_fd_sc_hd__a22o_1
X_1367_ net118 _0729_ _0730_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__and3_1
X_1298_ _0584_ _0216_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1797__220 vssd1 vssd1 vccd1 vccd1 _1797__220/HI net220 sky130_fd_sc_hd__conb_1
XFILLER_0_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput27 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xinput38 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1221_ team_11_WB.instance_to_wrap.sending.currentState\[3\] _0205_ _0206_ vssd1
+ vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__o21ai_1
X_1152_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[101\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[117\] vssd1 vssd1 vccd1
+ vccd1 _0695_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1083_ net346 net111 _0660_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0936_ team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[2\] _0474_
+ _0478_ _0580_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0867_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[15\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[14\]
+ team_11_WB.instance_to_wrap.sending.cnt_20ms\[16\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_24_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0798_ net315 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[0\] vssd1 vssd1 vccd1
+ vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1419_ net302 _0556_ net180 _0362_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_39_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1364__B1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 team_11_WB.instance_to_wrap.kp.buffertop.nrst vssd1 vssd1 vccd1 vccd1 net160
+ sky130_fd_sc_hd__buf_2
Xfanout171 net176 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_4
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1770_ net197 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XANTENNA__1726__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1769__196 vssd1 vssd1 vccd1 vccd1 _1769__196/HI net196 sky130_fd_sc_hd__conb_1
X_1204_ _0548_ _0554_ _0555_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__or4b_1
X_1135_ net383 net103 _0686_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__o21a_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1066_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[58\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[74\] vssd1 vssd1 vccd1
+ vccd1 _0652_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0919_ _0572_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold5 team_11_WB.instance_to_wrap.kp.controlstop.upper vssd1 vssd1 vccd1 vccd1 net265
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1822_ net153 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1753_ net248 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_53_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1684_ clknet_leaf_4_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keyvalid
+ net161 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.debouncertop.keyvalid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout175_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1118_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[84\] net137 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[100\] vssd1 vssd1 vccd1
+ vccd1 _0678_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1049_ net379 net103 _0643_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1817__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout88_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1805_ net225 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_14_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1736_ clknet_leaf_21_wb_clk_i _0192_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1667_ clknet_leaf_20_wb_clk_i _0177_ _0018_ vssd1 vssd1 vccd1 vccd1 team_11_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1598_ clknet_leaf_19_wb_clk_i _0112_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input20_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1521_ clknet_leaf_8_wb_clk_i _0035_ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[21\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1452_ net94 _0212_ _0335_ _0351_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[91\]
+ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__a32o_1
X_1383_ net54 _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1482__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1719_ clknet_leaf_12_wb_clk_i _0012_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1473__A2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0952_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\] net110 net85
+ _0594_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0883_ net117 _0544_ _0545_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1504_ net4 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1435_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[50\] _0339_ _0345_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[66\] _0376_ vssd1 vssd1
+ vccd1 vccd1 _0377_ sky130_fd_sc_hd__a221o_1
X_1366_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[15\] _0583_ _0264_
+ _0315_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__a31o_1
X_1297_ _0252_ _0253_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__or2_1
XANTENNA__1455__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_1_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1446__A2 _0341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput28 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput39 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1220_ team_11_WB.instance_to_wrap.sending.currentState\[3\] _0205_ vssd1 vssd1 vccd1
+ vccd1 _0207_ sky130_fd_sc_hd__nor2_1
X_1151_ net400 net103 _0694_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__o21a_1
X_1082_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[66\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[82\] net99 vssd1 vssd1
+ vccd1 vccd1 _0660_ sky130_fd_sc_hd__a221o_1
XANTENNA__1437__A2 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0935_ team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[1\] _0461_
+ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0866_ net309 _0531_ _0530_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[29\]
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0797_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[0\] _0491_ vssd1 vssd1 vccd1
+ vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[0\] sky130_fd_sc_hd__and2b_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1418_ _0357_ _0358_ _0359_ _0361_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1349_ _0296_ _0300_ _0301_ _0302_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_39_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1428__A2 _0342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout172 net173 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_2
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1419__A2 _0556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1203_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[9\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[11\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__and4b_1
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1134_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[92\] net137 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[108\] net95 vssd1 vssd1
+ vccd1 vccd1 _0686_ sky130_fd_sc_hd__a221o_1
X_1065_ net398 net103 net82 _0651_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout120_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0918_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\] _0551_ _0563_ vssd1 vssd1
+ vccd1 vccd1 _0572_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0849_ net312 _0522_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[21\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1337__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1224__S net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 net49 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1821_ net155 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1752_ net247 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_53_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1683_ clknet_leaf_0_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[7\]
+ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ net402 net113 _0677_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_0_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1048_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[49\] net144 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[65\] net95 vssd1 vssd1
+ vccd1 vccd1 _0643_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1688__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1833__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1761__256 vssd1 vssd1 vccd1 vccd1 net256 _1761__256/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_27_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1494__B1 _0345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1804_ net224 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1710__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1735_ clknet_leaf_10_wb_clk_i _0191_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1666_ clknet_leaf_10_wb_clk_i _0176_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1597_ clknet_leaf_21_wb_clk_i _0111_ net172 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1485__B1 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1828__A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input13_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1520_ clknet_leaf_25_wb_clk_i _0034_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1451_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\] _0346_ _0352_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[115\] _0384_ vssd1 vssd1
+ vccd1 vccd1 _0392_ sky130_fd_sc_hd__a221o_1
X_1382_ net55 net56 _0328_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1467__B1 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1718_ clknet_leaf_10_wb_clk_i _0011_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1649_ clknet_leaf_11_wb_clk_i _0159_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input5_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1458__B1 _0348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1449__B1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0951_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[1\] net145 net128
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[17\] vssd1 vssd1 vccd1
+ vccd1 _0594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0882_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[1\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[0\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _0545_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1503_ net3 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[6\]
+ sky130_fd_sc_hd__clkbuf_1
X_1434_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[10\] _0346_ _0349_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[18\] vssd1 vssd1 vccd1
+ vccd1 _0376_ sky130_fd_sc_hd__a22o_1
X_1365_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[7\] net90 vssd1 vssd1
+ vccd1 vccd1 _0315_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1296_ _0457_ _0240_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout150_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1128__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput29 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1150_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[100\] net137 net121
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[116\] net95 vssd1 vssd1
+ vccd1 vccd1 _0694_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1081_ net396 net109 _0659_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0934_ team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[2\] _0460_
+ _0478_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0865_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[27\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[26\]
+ _0442_ _0527_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0796_ _0481_ _0482_ _0487_ _0490_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__or4_4
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1417_ _0557_ _0356_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__or3_1
X_1348_ _0256_ _0278_ _0281_ _0238_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_39_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1279_ net264 _0236_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1836__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout140 net143 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout173 net176 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_4
Xfanout151 _0585_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1202_ _0722_ _0723_ _0720_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1133_ net391 net115 _0685_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__o21a_1
X_1064_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[57\] net144 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[73\] vssd1 vssd1 vccd1
+ vccd1 _0651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0917_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[9\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _0571_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0848_ _0521_ _0522_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[20\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0779_ _0476_ _0477_ _0478_ _0461_ net332 vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a32o_1
X_1787__210 vssd1 vssd1 vccd1 vccd1 _1787__210/HI net210 sky130_fd_sc_hd__conb_1
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7 net46 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1820_ net153 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1751_ net246 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_25_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1682_ clknet_leaf_0_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[6\]
+ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1500__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1116_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[83\] net149 net131
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[99\] net98 vssd1 vssd1
+ vccd1 vccd1 _0677_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1047_ net349 net107 net83 _0642_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1657__RESET_B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1803_ team_11_WB.instance_to_wrap.kp.controlstop.msg_tx_ctrl vssd1 vssd1 vccd1 vccd1
+ net52 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1734_ clknet_leaf_4_wb_clk_i _0190_ net161 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
X_1665_ clknet_leaf_10_wb_clk_i _0175_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1596_ clknet_leaf_24_wb_clk_i _0110_ net171 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout180_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1485__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1832__236 vssd1 vssd1 vccd1 vccd1 _1832__236/HI net236 sky130_fd_sc_hd__conb_1
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1508__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1450_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[27\] _0347_ _0389_
+ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__a211o_1
X_1381_ net56 _0328_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1717_ clknet_leaf_10_wb_clk_i _0010_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1648_ clknet_leaf_1_wb_clk_i _0158_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.controlstop.upper
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1579_ clknet_leaf_17_wb_clk_i _0093_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1672__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0950_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[8\] net107 net83
+ _0593_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1774__201 vssd1 vssd1 vccd1 vccd1 _1774__201/HI net201 sky130_fd_sc_hd__conb_1
XANTENNA__1082__C1 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0881_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[1\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[0\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _0544_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1502_ net2 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1433_ _0324_ _0363_ _0373_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__or4_1
X_1364_ _0308_ _0314_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[6\]
+ _0264_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__o2bb2a_1
X_1295_ _0457_ _0237_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_46_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout143_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_12_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1080_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[65\] net144 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[81\] net99 vssd1 vssd1
+ vccd1 vccd1 _0659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1523__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0933_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[13\] _0579_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.lcd_en sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0864_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[27\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[26\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[28\] _0527_ _0442_ vssd1 vssd1 vccd1
+ vccd1 _0530_ sky130_fd_sc_hd__a41o_1
X_0795_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[8\] _0488_ _0489_ vssd1 vssd1
+ vccd1 vccd1 _0490_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1416_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[8\] _0346_ _0352_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[112\] _0337_ vssd1 vssd1
+ vccd1 vccd1 _0360_ sky130_fd_sc_hd__a221o_1
X_1347_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\] net152 _0246_
+ _0441_ _0252_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1278_ net271 _0234_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_50_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout130 net134 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout174 net175 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_4
Xfanout152 _0583_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
Xfanout141 net143 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_2
Xfanout163 net166 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_4
Xfanout185 team_11_WB.instance_to_wrap.kp.buffertop.nrst vssd1 vssd1 vccd1 vccd1 net185
+ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1201_ _0717_ _0721_ team_11_WB.instance_to_wrap.sending.currentState\[5\] vssd1
+ vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1132_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[91\] net150 net133
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[107\] net98 vssd1 vssd1
+ vccd1 vccd1 _0685_ sky130_fd_sc_hd__a221o_1
X_1063_ net350 net107 net83 _0650_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__o22a_1
XANTENNA__1704__RESET_B net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0916_ _0569_ _0570_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0847_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[15\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[20\]
+ _0510_ _0519_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0778_ _0479_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout106_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 net43 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input36_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1750_ net245 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1681_ clknet_leaf_0_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[5\]
+ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1115_ net345 net112 _0676_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_0_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1046_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[48\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[64\] vssd1 vssd1 vccd1
+ vccd1 _0642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1697__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1494__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1802_ team_11_WB.instance_to_wrap.sending.lcd_en vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1733_ clknet_leaf_0_wb_clk_i _0189_ net156 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1664_ clknet_leaf_7_wb_clk_i _0174_ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1595_ clknet_leaf_23_wb_clk_i _0109_ net169 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout173_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1485__A2 _0346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1029_ net373 net104 _0633_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout86_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ team_11_WB.instance_to_wrap.kp.keypadtop.next_keyvalid _0491_ vssd1 vssd1
+ vccd1 vccd1 _0328_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1467__A2 _0336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0978__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1716_ clknet_leaf_10_wb_clk_i _0009_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1751__246 vssd1 vssd1 vccd1 vccd1 net246 _1751__246/LO sky130_fd_sc_hd__conb_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1647_ clknet_leaf_27_wb_clk_i _0157_ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1578_ clknet_leaf_13_wb_clk_i _0092_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1458__A2 _0345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1091__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1449__A2 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0880_ net117 _0542_ _0543_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1501_ net1 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[4\]
+ sky130_fd_sc_hd__clkbuf_1
X_1432_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[2\] _0340_ _0341_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[122\] vssd1 vssd1 vccd1
+ vccd1 _0374_ sky130_fd_sc_hd__a22o_1
X_1363_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\] net152 _0259_
+ net188 _0591_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a221oi_1
X_1294_ _0250_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_61_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ _0571_ _0578_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[11\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__a211o_1
X_0863_ net309 _0529_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[28\]
+ sky130_fd_sc_hd__xor2_1
X_0794_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[11\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[13\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[12\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__or4b_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1415_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[40\] _0336_ _0349_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[16\] _0355_ vssd1 vssd1
+ vccd1 vccd1 _0359_ sky130_fd_sc_hd__a221o_1
X_1346_ _0239_ _0243_ net187 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__o21a_1
X_1277_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[16\] _0234_ vssd1 vssd1 vccd1
+ vccd1 _0236_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1757__252 vssd1 vssd1 vccd1 vccd1 net252 _1757__252/LO sky130_fd_sc_hd__conb_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout120 net126 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout131 net133 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
Xfanout153 net155 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
Xfanout164 net166 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
Xfanout186 _0461_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_17_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1200_ _0717_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1131_ net370 net112 net86 _0684_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__o22a_1
X_1062_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[56\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[72\] vssd1 vssd1 vccd1
+ vccd1 _0650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0915_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[10\] _0567_ _0558_ vssd1 vssd1
+ vccd1 vccd1 _0570_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0846_ net318 _0520_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0777_ _0475_ _0477_ _0478_ _0463_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1329_ _0241_ _0238_ _0278_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold9 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[6\] vssd1 vssd1 vccd1 vccd1
+ net269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0942__A team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1680_ clknet_leaf_0_wb_clk_i team_11_WB.instance_to_wrap.kp.keypadtop.next_keycode\[4\]
+ net157 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1497__B1 _0349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1114_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[82\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[98\] net99 vssd1 vssd1
+ vccd1 vccd1 _0676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1045_ net351 net104 _0641_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1421__B1 _0338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0829_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[13\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[12\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[14\] _0506_ vssd1 vssd1 vccd1 vccd1
+ _0510_ sky130_fd_sc_hd__and4_2
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1412__B1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1479__B1 _0349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1801_ net223 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1732_ clknet_leaf_4_wb_clk_i _0188_ net161 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1663_ clknet_leaf_7_wb_clk_i _0173_ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1594_ clknet_leaf_13_wb_clk_i _0108_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout166_A team_11_WB.instance_to_wrap.kp.buffertop.nrst vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_1028_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[39\] net138 net122
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[55\] net97 vssd1 vssd1
+ vccd1 vccd1 _0633_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_24_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0757__A team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_1765__192 vssd1 vssd1 vccd1 vccd1 _1765__192/HI net192 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_34_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1164__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1809__229 vssd1 vssd1 vccd1 vccd1 _1809__229/HI net229 sky130_fd_sc_hd__conb_1
XANTENNA__1588__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1715_ clknet_leaf_10_wb_clk_i _0003_ net179 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1646_ clknet_leaf_27_wb_clk_i _0156_ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1577_ clknet_leaf_9_wb_clk_i _0091_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[77\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_64_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input11_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1500_ net266 net135 _0436_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1431_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[42\] _0336_ _0348_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[74\] vssd1 vssd1 vccd1
+ vccd1 _0373_ sky130_fd_sc_hd__a22o_1
XANTENNA__1137__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1362_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[5\] net90 _0308_
+ _0313_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__a22o_1
X_1293_ _0020_ _0021_ _0001_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout129_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1629_ clknet_leaf_25_wb_clk_i _0001_ net158 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input3_A gpio_in[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0931_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[5\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[4\]
+ team_11_WB.instance_to_wrap.sending.cnt_500hz\[7\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_31_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0862_ _0528_ _0529_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[27\]
+ sky130_fd_sc_hd__nor2_1
X_0793_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[14\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[17\]
+ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_21_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1414_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[120\] _0341_ _0347_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[24\] _0354_ vssd1 vssd1
+ vccd1 vccd1 _0358_ sky130_fd_sc_hd__a221o_1
X_1345_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[2\] _0299_ _0264_
+ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1276_ _0234_ _0235_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0740__D net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout121 net126 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_2
Xfanout110 net116 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_2
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout143 net151 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
Xfanout176 net185 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
Xfanout187 team_11_WB.instance_to_wrap.kp.controlstop.mode vssd1 vssd1 vccd1 vccd1
+ net187 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1130_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[90\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[106\] vssd1 vssd1 vccd1
+ vccd1 _0684_ sky130_fd_sc_hd__a22o_1
X_1061_ net341 net110 _0649_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0914_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[10\] _0567_ vssd1 vssd1 vccd1
+ vccd1 _0569_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0845_ net300 _0520_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[19\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1713__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0776_ team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[0\] _0472_
+ _0473_ net186 vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1328_ _0459_ _0001_ _0020_ _0261_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__o31ai_2
X_1259_ net290 _0224_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1794__217 vssd1 vssd1 vccd1 vccd1 _1794__217/HI net217 sky130_fd_sc_hd__conb_1
XFILLER_0_62_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1113_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[89\] net109 net85
+ _0675_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_49_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1044_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[47\] net145 net122
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[63\] net96 vssd1 vssd1
+ vccd1 vccd1 _0641_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0828_ net301 _0508_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[13\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0759_ team_11_WB.instance_to_wrap.kp.debouncertop.next_receive_ready team_11_WB.instance_to_wrap.kp.debouncertop.receive_ready
+ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0999__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input41_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1800_ team_11_WB.instance_to_wrap.sending.lcd_rs vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1731_ clknet_leaf_4_wb_clk_i _0187_ net161 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_2
X_1662_ clknet_leaf_7_wb_clk_i _0172_ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1593_ clknet_leaf_9_wb_clk_i _0107_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[93\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1027_ net401 net113 net87 _0632_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout159_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1149__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[64\] vssd1 vssd1
+ vccd1 vccd1 net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1714_ clknet_leaf_3_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[29\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1645_ clknet_leaf_1_wb_clk_i _0155_ net157 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1576_ clknet_leaf_26_wb_clk_i _0090_ net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1430_ net268 net135 net168 _0372_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__o211a_1
X_1361_ _0259_ _0309_ _0310_ _0312_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__a31o_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
X_1292_ net187 _0590_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1628_ clknet_leaf_27_wb_clk_i _0000_ net160 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1559_ clknet_leaf_18_wb_clk_i _0073_ net174 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0930_ net339 net38 net40 vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__and3b_1
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0861_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[27\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[26\]
+ _0527_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0792_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[1\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[0\]
+ _0485_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1413_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[0\] _0340_ _0344_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[80\] _0353_ vssd1 vssd1
+ vccd1 vccd1 _0357_ sky130_fd_sc_hd__a221o_1
X_1344_ _0261_ _0282_ _0295_ _0298_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__o22a_1
X_1275_ net285 _0232_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout141_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1451__C1 _0384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout122 net126 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout111 net116 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
Xfanout100 _0589_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_2
Xfanout155 net76 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout144 net145 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
Xfanout133 net134 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_2
Xfanout188 team_11_WB.instance_to_wrap.kp.controlstop.mode vssd1 vssd1 vccd1 vccd1
+ net188 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout166 team_11_WB.instance_to_wrap.kp.buffertop.nrst vssd1 vssd1 vccd1 vccd1 net166
+ sky130_fd_sc_hd__buf_2
Xfanout177 net185 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1060_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[55\] net145 net128
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[71\] net98 vssd1 vssd1
+ vccd1 vccd1 _0649_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0913_ _0567_ _0568_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__nor2_1
X_0844_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[15\] _0510_ _0519_ vssd1 vssd1
+ vccd1 vccd1 _0520_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0775_ team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[2\] _0472_
+ _0473_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1327_ _0250_ _0281_ _0256_ _0441_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__a211oi_1
X_1258_ _0224_ _0225_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__and2_1
X_1189_ net295 net96 _0713_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1430__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1497__A2 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1747__242 vssd1 vssd1 vccd1 vccd1 net242 _1747__242/LO sky130_fd_sc_hd__conb_1
XFILLER_0_45_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1112_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[81\] net144 net127
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[97\] vssd1 vssd1 vccd1
+ vccd1 _0675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1043_ net406 net114 net87 _0640_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_29_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1421__A2 _0336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ _0508_ _0509_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[12\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout104_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0758_ team_11_WB.instance_to_wrap.kp.debouncertop.next_receive_ready team_11_WB.instance_to_wrap.kp.debouncertop.receive_ready
+ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__and2b_2
XFILLER_0_40_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1488__A2 _0556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1412__A2 _0342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1604__RESET_B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input34_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1479__A2 _0348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1818__232 vssd1 vssd1 vccd1 vccd1 _1818__232/HI net232 sky130_fd_sc_hd__conb_1
XFILLER_0_26_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1730_ clknet_leaf_12_wb_clk_i _0186_ net180 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.lcd_rs
+ sky130_fd_sc_hd__dfrtp_1
X_1661_ clknet_leaf_7_wb_clk_i _0171_ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592_ clknet_leaf_22_wb_clk_i _0106_ net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1026_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[38\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[54\] vssd1 vssd1 vccd1
+ vccd1 _0632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1330__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold91 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[55\] vssd1 vssd1
+ vccd1 vccd1 net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[16\] vssd1 vssd1
+ vccd1 vccd1 net340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1526__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1713_ clknet_leaf_3_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[28\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1644_ clknet_leaf_0_wb_clk_i _0154_ net157 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1575_ clknet_leaf_18_wb_clk_i _0089_ net176 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout171_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1009_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[37\] net106 net91
+ _0623_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout84_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
X_1360_ team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl _0590_ _0260_
+ _0311_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a211o_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
X_1291_ _0001_ _0021_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1707__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1627_ clknet_leaf_24_wb_clk_i _0141_ net159 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_1558_ clknet_leaf_20_wb_clk_i _0072_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_1489_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[127\] _0341_ vssd1
+ vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1460__B1 _0347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0860_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[26\] _0527_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[27\]
+ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0791_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[4\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[6\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[5\] vssd1 vssd1 vccd1 vccd1 _0486_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_3_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1412_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[32\] _0342_ _0350_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[56\] vssd1 vssd1 vccd1
+ vccd1 _0356_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1343_ _0296_ _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__or2_1
X_1274_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[15\] _0232_ vssd1 vssd1 vccd1
+ vccd1 _0234_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1451__B1 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0989_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[27\] net112 net85
+ _0613_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout112 net116 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_2
Xfanout101 net108 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_4
Xfanout134 _0586_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_2
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net151 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_2
Xfanout167 net169 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
Xfanout178 net185 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1629__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0912_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[9\] _0566_ _0558_ vssd1 vssd1
+ vccd1 vccd1 _0568_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0843_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[17\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[16\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[19\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0774_ team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[1\] _0474_
+ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1326_ _0250_ _0281_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__and2_1
X_1257_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[7\] _0223_ vssd1 vssd1 vccd1
+ vccd1 _0225_ sky130_fd_sc_hd__or2_1
XANTENNA__1722__RESET_B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1188_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[119\] _0460_ net139
+ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1424__B1 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1415__B1 _0349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1111_ net359 net105 net83 _0674_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1042_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[46\] net148 net132
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[62\] vssd1 vssd1 vccd1
+ vccd1 _0640_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0826_ net324 _0506_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0757_ team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl vssd1 vssd1 vccd1
+ vccd1 _0459_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1309_ _0441_ _0590_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1660_ clknet_leaf_6_wb_clk_i _0170_ net165 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.sending.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1591_ clknet_leaf_18_wb_clk_i _0105_ net176 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1784__207 vssd1 vssd1 vccd1 vccd1 _1784__207/HI net207 sky130_fd_sc_hd__conb_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1025_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[45\] net106 net91
+ _0631_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0809_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[4\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[5\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[6\] _0494_ vssd1 vssd1 vccd1 vccd1
+ _0498_ sky130_fd_sc_hd__and4_1
X_1789_ net212 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_4_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1772__199 vssd1 vssd1 vccd1 vccd1 _1772__199/HI net199 sky130_fd_sc_hd__conb_1
XFILLER_0_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold70 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[16\] vssd1 vssd1 vccd1 vccd1
+ net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[63\] vssd1 vssd1
+ vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[86\] vssd1 vssd1
+ vccd1 vccd1 net352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1712_ clknet_leaf_3_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[27\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1566__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1643_ clknet_leaf_0_wb_clk_i _0153_ net157 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1574_ clknet_leaf_20_wb_clk_i _0088_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout164_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1008_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[29\] net141 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[45\] vssd1 vssd1 vccd1
+ vccd1 _0623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
X_1290_ _0245_ _0246_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1626_ clknet_leaf_14_wb_clk_i _0140_ net183 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_1557_ clknet_leaf_22_wb_clk_i _0071_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_1488_ net382 _0556_ net182 _0425_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_0__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_53_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0790_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[3\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[2\]
+ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[7\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1411_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[64\] _0345_ _0351_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[88\] vssd1 vssd1 vccd1
+ vccd1 _0355_ sky130_fd_sc_hd__a22o_1
X_1342_ _0238_ _0252_ _0281_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__mux2_1
X_1273_ _0232_ net278 vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1451__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout127_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0988_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[19\] net147 net130
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[35\] vssd1 vssd1 vccd1
+ vccd1 _0613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout102 net108 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout113 net115 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_2
X_1609_ clknet_leaf_10_wb_clk_i _0123_ net178 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[109\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout135 _0556_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_4
Xfanout146 net151 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
Xfanout124 net126 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
Xfanout179 net181 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_4
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_4
Xfanout157 net160 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input1_A gpio_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1669__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0911_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[8\] team_11_WB.instance_to_wrap.sending.cnt_500hz\[9\]
+ _0563_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__and3_1
X_0842_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[18\] _0517_ net299 vssd1 vssd1
+ vccd1 vccd1 _0518_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0773_ team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[1\] _0472_
+ _0473_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1325_ _0001_ _0020_ _0021_ net188 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1256_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[7\] _0223_ vssd1 vssd1 vccd1
+ vccd1 _0224_ sky130_fd_sc_hd__nand2_1
X_1187_ net317 net115 net88 _0712_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1110_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[80\] net140 net124
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[96\] vssd1 vssd1 vccd1
+ vccd1 _0674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1041_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[53\] net106 net91
+ _0639_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0825_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[12\] _0506_ vssd1 vssd1 vccd1
+ vccd1 _0508_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0756_ _0457_ _0458_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl
+ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1308_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[0\] net90 vssd1 vssd1
+ vccd1 vccd1 _0265_ sky130_fd_sc_hd__nand2b_1
X_1239_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[7\] net283 net186 vssd1
+ vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1777__204 vssd1 vssd1 vccd1 vccd1 _1777__204/HI net204 sky130_fd_sc_hd__conb_1
XFILLER_0_38_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1590_ clknet_leaf_19_wb_clk_i _0104_ net173 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1024_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[37\] net141 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[53\] vssd1 vssd1 vccd1
+ vccd1 _0631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0808_ _0491_ _0496_ _0497_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[5\]
+ sky130_fd_sc_hd__and3_1
X_1788_ net211 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
X_0739_ net5 vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold60 team_11_WB.instance_to_wrap.sending.cnt_20ms\[3\] vssd1 vssd1 vccd1 vccd1
+ net320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[76\] vssd1 vssd1
+ vccd1 vccd1 net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[18\] vssd1 vssd1
+ vccd1 vccd1 net331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[17\] vssd1 vssd1
+ vccd1 vccd1 net353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1711_ clknet_leaf_3_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[26\]
+ net164 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1642_ clknet_leaf_0_wb_clk_i _0152_ net157 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1573_ clknet_leaf_21_wb_clk_i _0087_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_1007_ net348 net101 _0622_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout157_A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__clkbuf_4
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1625_ clknet_leaf_9_wb_clk_i _0139_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[125\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1556_ clknet_leaf_15_wb_clk_i _0070_ net178 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_1487_ _0419_ _0421_ _0422_ _0424_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_53_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1460__A2 _0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[48\] _0339_ _0348_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[72\] vssd1 vssd1 vccd1
+ vccd1 _0354_ sky130_fd_sc_hd__a22o_1
X_1341_ net188 _0250_ _0253_ _0284_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__a31o_1
X_1272_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[13\] _0230_ net277 vssd1 vssd1
+ vccd1 vccd1 _0233_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1451__A2 _0346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0987_ net369 net109 net85 _0612_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1550__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1608_ clknet_leaf_22_wb_clk_i _0122_ net168 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0962__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout103 net108 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__buf_2
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout136 net139 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_2
X_1539_ clknet_leaf_24_wb_clk_i _0053_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[39\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout147 net151 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_2
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
Xfanout114 net115 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_2
Xfanout169 net176 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
Xfanout158 net160 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_4
X_1805__225 vssd1 vssd1 vccd1 vccd1 _1805__225/HI net225 sky130_fd_sc_hd__conb_1
XFILLER_0_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0953__A1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0910_ _0566_ net117 _0565_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__and3b_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0841_ net297 _0517_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[18\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0772_ _0472_ _0473_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1324_ _0242_ _0257_ _0276_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__o21ba_1
X_1255_ _0443_ _0222_ _0223_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1186_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[118\] net148 vssd1
+ vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1424__A2 _0340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1360__A1 team_11_WB.instance_to_wrap.kp.controlstop.next_msg_tx_ctrl vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1415__A2 _0336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1040_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[45\] net141 net123
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[61\] vssd1 vssd1 vccd1
+ vccd1 _0639_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1754__249 vssd1 vssd1 vccd1 vccd1 net249 _1754__249/LO sky130_fd_sc_hd__conb_1
X_0824_ _0506_ _0507_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[11\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0755_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[1\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[0\]
+ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[2\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__or4b_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1307_ _0263_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__inv_2
X_1238_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[6\] net293 net186 vssd1
+ vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1169_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[117\] net107 net92
+ _0703_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1653__RESET_B net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1023_ net361 net101 net82 _0630_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_wb_clk_i clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1787_ net210 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0807_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[4\] _0494_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__a21o_1
X_0738_ team_11_WB.instance_to_wrap.sending.cnt_500hz\[3\] vssd1 vssd1 vccd1 vccd1
+ _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout102_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input32_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[25\] vssd1 vssd1 vccd1 vccd1
+ net310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[4\] vssd1 vssd1 vccd1
+ vccd1 net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 team_11_WB.instance_to_wrap.kp.controlstop.previous_key_count\[0\] vssd1 vssd1
+ vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 net53 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[22\] vssd1 vssd1
+ vccd1 vccd1 net354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1490__B1 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1790__213 vssd1 vssd1 vccd1 vccd1 _1790__213/HI net213 sky130_fd_sc_hd__conb_1
X_1710_ clknet_leaf_3_wb_clk_i team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[25\]
+ net162 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.count\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_1641_ clknet_leaf_0_wb_clk_i _0151_ net156 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1572_ clknet_leaf_9_wb_clk_i _0086_ net177 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1575__RESET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1006_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[28\] net136 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[44\] net95 vssd1 vssd1
+ vccd1 vccd1 _0622_ sky130_fd_sc_hd__a221o_1
XANTENNA__1481__B1 _0345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1839_ net238 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_0_60_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1472__B1 _0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1553__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__clkbuf_4
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1463__B1 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1624_ clknet_leaf_23_wb_clk_i _0138_ net167 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1555_ clknet_leaf_16_wb_clk_i _0069_ net170 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1486_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[102\] _0343_ _0350_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[62\] _0423_ vssd1 vssd1
+ vccd1 vccd1 _0424_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1762__189 vssd1 vssd1 vccd1 vccd1 _1762__189/HI net189 sky130_fd_sc_hd__conb_1
XFILLER_0_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout82_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1445__B1 _0344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1340_ _0243_ _0277_ _0278_ _0255_ _0294_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_20_wb_clk_i clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_1271_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[13\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[14\]
+ _0230_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1436__B1 _0351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0986_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[18\] net146 net129
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[34\] vssd1 vssd1 vccd1
+ vccd1 _0612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1607_ clknet_leaf_17_wb_clk_i _0121_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout104 net108 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_2
Xfanout126 _0586_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_2
XANTENNA__1590__RESET_B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 net139 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xfanout115 net116 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_2
X_1538_ clknet_leaf_14_wb_clk_i _0052_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[38\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_4
X_1469_ _0210_ _0317_ _0340_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__a2bb2o_1
Xfanout148 net150 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_38_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1427__B1 _0352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0840_ _0516_ _0517_ vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.clkdivtop.next_count\[17\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0771_ _0464_ _0467_ _0468_ _0469_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_58_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1323_ _0001_ _0021_ _0246_ net188 vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__o211a_1
X_1254_ team_11_WB.instance_to_wrap.sending.cnt_20ms\[5\] team_11_WB.instance_to_wrap.sending.cnt_20ms\[4\]
+ team_11_WB.instance_to_wrap.sending.cnt_20ms\[6\] _0538_ vssd1 vssd1 vccd1 vccd1
+ _0223_ sky130_fd_sc_hd__and4_1
X_1185_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[125\] net107 net92
+ _0711_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1409__B1 _0343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0969_ net353 net104 _0603_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1700__RESET_B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1768__195 vssd1 vssd1 vccd1 vccd1 _1768__195/HI net195 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_2_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0823_ net308 _0504_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0754_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[5\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[4\]
+ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[6\] team_11_WB.instance_to_wrap.kp.buffertop.keycode\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__or4b_4
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1306_ _0441_ _0247_ _0250_ _0262_ _0460_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1237_ team_11_WB.instance_to_wrap.kp.buffertop.keycode\[5\] net292 net186 vssd1
+ vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1168_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[109\] net142 net125
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[125\] vssd1 vssd1 vccd1
+ vccd1 _0703_ sky130_fd_sc_hd__a22o_1
X_1099_ net335 net111 _0668_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1693__RESET_B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1022_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[36\] net136 net119
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[52\] vssd1 vssd1 vccd1
+ vccd1 _0630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1786_ net209 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_0806_ team_11_WB.instance_to_wrap.kp.clkdivtop.count\[4\] team_11_WB.instance_to_wrap.kp.clkdivtop.count\[5\]
+ _0494_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__nand3_1
XFILLER_0_40_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0737_ net333 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1513__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 _0518_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 team_11_WB.instance_to_wrap.sending.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ net333 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold51 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[123\] vssd1 vssd1
+ vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[120\] vssd1 vssd1
+ vccd1 vccd1 net322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[113\] vssd1 vssd1
+ vccd1 vccd1 net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[19\] vssd1 vssd1
+ vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1640_ clknet_leaf_1_wb_clk_i net287 net157 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.buffertop.keycode_previous\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1571_ clknet_leaf_17_wb_clk_i _0085_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1005_ net374 net112 _0621_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1544__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1838_ net154 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1769_ net196 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1623_ clknet_leaf_17_wb_clk_i _0137_ net175 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1554_ clknet_leaf_14_wb_clk_i _0068_ net182 vssd1 vssd1 vccd1 vccd1 team_11_WB.instance_to_wrap.kp.decodertop.data_received\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1485_ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[14\] _0346_ _0352_
+ team_11_WB.instance_to_wrap.kp.decodertop.data_received\[118\] _0319_ vssd1 vssd1
+ vccd1 vccd1 _0423_ sky130_fd_sc_hd__a221o_1
.ends

