/*
* This is a template for your top level test bench!
* You are responsible for having a test bench for your top
* level design. Otherwise, your design will not be part
* of the tape-out.
*
* Please also include test benches for your team_02_WB
* and team_02_Wrapper modules, if needed to verify
* interfacing with the Wishbone Bus.
*
* The command to run this test bench is:
* make tbsim-source-team_02-team_02
*/

`timescale 1 ns / 1 ps

module team_02_tb();

    ///////////////////////////////////
    // Write your test bench code here!
    ///////////////////////////////////

endmodule